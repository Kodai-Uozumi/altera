��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���a?K���J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-@���rahZ����*��/}{�_@1������{S�������<�w$ɨ�h���G�m6
�DR���8�+I�S��n�D�N�����N�8t�>�Hc;��|B|X����}��_��t�ս߸�Z�C	�a1ﲀZ���dJh2-jwG�CUG@�t�k�k'v��ǔ{�q�%O���t����t�D�~w����+�#���]�0��mS��m%B����Ӻ��,Q�Q�?uG�Qy�����Q�Y�Bݣٳ���� [��(�� %����
�?<�곦���q1��B�ceH��.���s6�kk�`��y��&������i��0+�M��L,��.K��C���@J{�"F�6r/	�Y�B!zZ��۸9ߤ�Ha���3����!�L���!�`�(i3!�`�(i3���ue���!�`�(i3!�`�(i3F^I�i<}�sȸ�"rR!�`�(i3�4&8��z�[�X��ņ�3\SrXtN����f�%;.�J}��Ut���c�&��j�b�,t,�y�WW�W�ck��=~Ì��O�K�"��)�1������1������R���l%�odYǭ�%�Z[K�1��������;I6l��7�GQ�C����5�sȸ�"rR�· ���4���w0�DT��b֤�]�G�6���7��$�7��$EԔ	�8��6?���W+X�~{˕vC�|�ˏ8[$0�I�'�z��9���
�n|s�)>��!��<�ڒ�]X/��~�5:��fĝke�!�`�(i3J��+GP��fhH�{V�RDFR7�?D��׊�'�t+��u��^�ץ�7z��	.�V�~�-���\�>�/E�CԵ�_�*���d��4D���t���װh����t�D�R�WZ��@O���t��A�Pf�d�:o+'�E}u1�R�Ȫ~���		�X.]���}�W��� ���G���p�@OM.Ir��"���tc��=�����?�o�JH�S�Zt�(���b?(���&�!+5���Y�҃ڹ�^��2���96v_ �7�����T�٥��T)'��:�Jl
��Pn�߶h��Myf%���G�v���Y�p+�~��]a�{��>LTd��e�R��b�7S�����i�F��2�+g�@7��cؖ�r�M�?��	4�����wƃ(%��<'����Z"}�p����>�UKW�*�	S&&�s m�Ht���11
����}C9�S�+o���oBg�Caz�~�?���Bꮷ����A?�>�Q�k^�Á�)�o��.&l��ʩ�R'���=�\�W�EC�)�6-��~h�ӦI%}���/�çEF�)�]ܤ�1�G�Qc}y�����߫��Ѷm��Ǹ�vJ]�3�<
d�>��W����`�r����Fz�NK8�y �����<7u!�`�(i3f�s�J!�`�(i3NK8�y ��K�"��)�ul֗��|�!�`�(i3!�`�(i31������!�`�(i3&��潹!�`�(i3m�7�TG���^:��lFE�߇ç�b� ��Jײ?����!�`�(i3�m��7E��!�`�(i3!�`�(i3?������ޝq�~�[_.H P긭so3#���^�_!��� ���r�>��f1~�?��Ӑ����~�f h,��3h!�`�(i3!�`�(i3�· ���4!�`�(i3��J���FB���Շd��@Ő��t勪�i�/��{�P:tg��ݖ˘�&��Lӳ��{%_��6�z�
^��t&�"��+E�Tw�· ���4!�`�(i3h,��3h!�`�(i3!�`�(i3�· ���4m6
�DR�П�� j�L*կ`��%�����-���,���x��
R���eU<�������|[���HHi���~����Us��9�ۗ�蠒pP��!�`�(i3!�`�(i31������!�`�(i3&��潹!�`�(i3�����,I��Y7h�dČ���4�B��ٴ��s±���w	Qrk)F9�>�^W+X�~{��2�N��T$q��mKx"E&��� ���yoZ�P/Y�l��aLR����|���\X�TQ���EW�)U���a���C��iF�9�����$���y�VJ!���(�a��ܡ\{S�@g�(4������j��Z&��Ûf��O�.��+Y�B�&�%u�<��6u�G	O�V�g���ޔ��(p�]�u��.tƲ����%���a�>��$d�I�v���v,���h���ur�}w�*W+X�~{�ւ���z�X,mvvԩ|PM��!����E:v��M��n���/刲�Z��Utu⯃�ic" le�j�@���p��}K��f<�,=K�F~�?|�[_X��ˆk�=c�!8�Ԏi��p�7��Z鎬������~/[�� &He�ߏ=W�֯�^��N�&��?�2�1p�Qk�� h��ߖ�g��o�4��?����DNZ�j׫���?_W�\I��ఽ��`g�5��!08�tw:g�/�6=m�	n� ^�d�#2��0�DQ�L���EuZoO�=����'�ނ�ebÆ���p��'��aC�h�>�4����CX36-Q��ܹ��E!����梡���h�3��3%��׍����}0�st&���\�vūx`��:�֡�\�<7�X�e���V!���IÙ=�H�l��3d�`.�/'�����W;5B5Y+� �i7�sp>��=D3�OO�@I�I�z%��;5B5Y+�T�����N��=D3�OO~G��;ؔ�V@��n����&��J�f����t�Xx�s]���uC#����
p��#�IÙ=�H�&8���l�mq���)�:��j8HQ��e�z���V�RDFR7������`��I�t?�_��B�e�D�*�Y�p�Yч���Ҟ�+���A��33�V���C��\����<�(p�M�=�U� ���_~�?���4�ͻs�	Õ�)X�JK�IE��q{�f��a�:&�>��sH�2Da���`�M7Э7l��A���ZL�4��L��Q<G�^���_%���}����Eڑi
�樄�ZWu)�=>�q�E#�U7�D�>���RQ�˕��~G��;ؔ��r�C©���+7IÙ=�H��`�Sb�j|~��A�!`�u�!j�4I^J<�
� �>׍�vA���P`�|��K�z��5��8�tʆ�In��t28�/�>��L�+�M�R��x���hA�q:i@_��R��w5�tF�~��j.o�c�\.U1+]�{r�J����{�OF8w�DƉqaݾ'���ߌ[����6�d�٣��c�A�L'b-a��K[.9�V���i|Stߛ�mBp�S��JHn��z��r9�3��\P�/vփZ���0�q{�f��a��{oS�6 �P�{0�7��65���5��8�t��\�v�I���#��������PPV��"tXۓښ-x�]�V����qG�d�w��V%�piS�G���HaM��-����׋4>&:��Op�M+�	�$<zL͊�q���b�Kzb���}g��u"��*�ΊJ~��ڹ 	��\�v��wc�}�![vl�+��3�-�#���[�3��z�/��;5B5Y+��\ԅ����i�@�t��c��1�u�K|]���TI�uK���j\C����)|fvl�+��3�-�#���[��0c(��<>p����ct�q�p�P���YG�zL͊�q�����������r���aM"��N�߄�4�X�)Х��؊�K�H��\�v��wc�}�![vl�+��3�-�#���[���d�%X!ԱX�|�O*)y
���z���n�؅��FJ��KL�IO�!ivl�+��3�-�#���[���)gΔc�G���`NOE���yn2�@F�4��d��X���n�R�[̈���d L��s�XS� �F�s��M_�_���wg�|��].��'���XwSn����P>7Xl����]�Jg����-c �ЄW:��2�-4�������A{��JVjN�h�Q�;������;��B�ip��{l�f|����%Hl�>���_�Z1~�g]�I���B��!nJ�Q�-Y���".7�!n}y���q���U��F�R�M�so�	�C�/ɽs���܉-`�6��+��us�Pc��?@W�m!��ʧ�9�x�^4/��?Ev�~������]�!��ѩ	 7l�"b��"am��%��{l�f|�ό���.Ӡ���f~��n��7�|��].��'���Xw�|���E�+kg�s��]b�|��].��'���Xw��]v�A�5P^�\8	���-�$�<��z��}�Q2�+�Yɶg�Y_���n��7�|��].��'���XwE�%5S��|���kJ�|��].��'���Xw��"N(�MO���t���x,pk�0��=��5t��vv�~������]�!��	Ǹ�y85��d!+��T��b�!cI��:F�X?�g��U-�eS2o�E�t��6�z�
^��̠ӷJė/�Ҏ��^�  @��:�2�{k�_V�\#V f�Lu�mE{le��K��ҋX����0�a1i~J����Ew(�9V(;�&����օP0��p�Q�@��߿�È�<�6&�nw���]�!�����#e��H^���P2<WV�㤚`3���j�ho���`-���z�f�Š,�%��p��qrۤG�#r�\���(.���*�KKZ鎬�������(����ｗ��u��;e5V�]C��( _�O
�_�Z)<��)�A�'z4ӭs��'K� Y�����r�_`��0#��=�8:~�� �d�OMb�O�Y�M�?�|��].��'���Xw�{ƕ��w���'�#&7Q�w�D�o��&Y��V��(��ug�X���K{��,cI��S}Ht�+37/�+�m�r�d ��(�
t�ژq���U����#��mW[�Ƶ\�rK�@<,у7G#+��Q2�+�Y�6UQ�㔩�S�(��ɒ���9�dMbZ鎬������fu��V�:Y3Iz�SŞ�Ӣ�8k>6s����]�!�����&��<o!f�	�Ĳb�M� �{�6�vg;Je'���Xw�j�7��o�${U��w�X�|0��X��������`y�����-x�~}0��/�0,�WT�j
�I��w��,c�A�L'� �3�,���BT�^��a(􆿳��[ihC�����։�s/�)���R8&���9�dMbZ鎬�������(���y�T�g}���`�L�iַ:���N3!�U\���<�����,�8��(�
t��Y�{'%s�h�v����}g��u"��*�ΊJ�˷���T�\ �ͪ�c�$�B"�c�z�
���8Z�6�vg;Je'���Xw���e�K�ѕ��J��<�..�4�ኈ�8���K(��z�j�;9�e��/}{�_@1�����&��H�˦�\��~T�����DM����p.s��|� �f׿���$	n��s�I�H/�v�6���l �;ۂ��IÙ=�H"�t�ѵ$r���@	Q�č�Y�����&��J�������׻P��#Y�dL�|�u0x�]�V��e�����1~��j.o�����i�]�!��	Ǹ�y85�>T
BFa@#e�����1~��j.o�c�\.U1+]d�TpubMpIÙ=�H���:ipSVUioέ���K�IE��;5B5Y+� �i7�sp>���=��s*c�r�w����bU^���j�b?u |�V���r�^�y4fCx=�a�ߩJ�9��č�Y���S�)37J*u�v3���?B]z�����B*�2���u���d��O�Z�:����!n�������s�3�t8��5���dq��}hU��xz��osq���{l�f|����%Hl�3�[i�`#��E<�J��yoZ�P/��A�,F��v_}���2
��;���GU���|kv�~������]�!�����#e��j�b��A�,�O
ɝe�{�f�U�V^q2��gͼs��Ę�}��U��Ÿ|��].��'���Xwu��:���hx��W����c��a�$Z%���*�k8���Hm�č�Y���S�)37J*u)T{6T'��ՁO�#d�č�Y���S�)37J*uc�A�L'��!�a�&H�[&-n�g��U-�e`�gB��,���Ξ1�R.%:7	v�.�f�3���u++J)tf��k�8�H3=-��7��B�>�9��(�
t�ژq���U��,���Ξd�$�j�|J�E�$tv�.�f�3�^-���Wm�_�����t���2E!^��@��1�@ �~)��*/�|�!���_- �v�j=U�h�]�vv���E�fZ@IE�U����S8��m�o�&i~G��;ؔa��-)�]��V+m�}.�Q�º�F����U�D�>i�ל�I�p\�WB����&�?T0�oKG�:nܑr�_@r�|S�Ǔ���aD�orǟD�uiL${?�����>��yܛ�	��|��	(���zL͊�q���19TH���'�3�$ �#^�Vn�^ֻ����XP��Ȼ4�t=�j�.�/'�����W;5B5Y+� �i7�sp>�
� �F״��`B캶S�)k��'n�^0o����SVc�Iۣ<�;�'��-d�Ryʆ�In��t�wc�}�![۟D�$0+�(ԛ���\�v��wc�}�![���z��>x��F�\.��0�q:i@_�8x<�A!tr��8`S�*���X���^ m�Z鎬�������(����5�	��]�k�K�ָ������Z�]�O�"�"m;��U6�k�#��.���t�:��F{iY;��'n�^0oޖW�/�
�^�=�Q�9�θ�c}k�,���Ξ1�R.%:7	v�.�f�3���u++J)t��V�b}1�MԲ����!n}y���q���U�S]�}�g��$y�z��eU�e�������&�Ժ����R
���rPޯ��-�0����'I']�5X�vZ��Bv�~������]�!�����#eH$�DZ� ��o30�@Cd�$�j����"�YVķ�;�����G�c�J�!�Ӑ��3�ql��J��{l�f|����%Hl��,���Ξd�$�j�|J�E�$tv�.�f�3��1h��*�1�צ�);[r�����R]Y�~�����ҋX���� 
���u���� �������9�O���Òx8�!��K��J<W�f�ӊ[�k碝{l�f|�ό���.�k:j%]a6��w%e���{l�f|��rs�i�jf� l�ǉ��F1x,0=]^	�&���Øf���t���2���B�|��m|�z��e�i�"�����{����c�Ļ�+�m�r�d ���9�dMbZ鎬��������E����X)���$U�����m|�Q'xF�#�
W/7�䬢�
���D/5xM�����?��9)J Ւ�&����i�{�#�	�����1p�Zc]�y���7G#+�Ǘ0z�cUL�n+q����`B�� {�>|wՓ8���/�H3�%9�5ܤ�@�@yo�8�@I}��A�"�b���"v�I��#��@f׿���$	n��s�xՉ�T�Ұ>D�c�lQKݗZ:���'n�^0o����y�]֡�\�<7�X�e���V!���IÙ=�H�]ƭ��&d&(C�#�7#^�Vn�^ֻ����XP���E)
i����$�b��ev�~�����M�-��#�Ay0Hb�Z'�2%;5B5Y+��q	k���A�O����!;�Y"f��g�o&�Y��>�_����6����?�y)��;ۂ���d�����#��QU(�M�z��K��J<W�f�ӊ[�k碝{l�f|�ό���.�k:j%]a6��w%e���{l�f|��rs�i�jf� l�ǉ��F1x,0=]^	�&������*��p��U�d�K��@�!n}y��Y�{'%s43u�R��}/A;T�c���Y#?M��^e@��V�m�C��x�T�\ ���p�N0��g��?`-ʂE�����7G#+�ǟ
��|�6|�+�� VU+I���(Bt|�x���� ��ѕ��J�� f�Lu�m�/
����X� L�u�۽t|Y�f�s�m��n��&�7a	��������W;5B5Y+� �i7�sp>��ߪ��ʙ��BC?T�<o�nïi�JHn��z��r9�3�ͫ��;���^hq��:�}0�st&���\�vūx`��:�7γҬ�,;r�mR-AFɈf�=K�:���A0���zk��p`V-u9�`�JHn��z��y`E���*`�"�X�� [3[��?;5B5Y+��4"�I<a�kGQ��l�4��H���^ֻ����XP����؇��7��'���ߌ[R)Ms	[����d���
zL͊�q��������Rm�Ƈ�hʨ}s����=Y��_�0z�cUL�ӒN��G�g�tNw��[
�}3���M:��2�8���Hm�č�Y���S�)37J*u��xc�lf#�}N9�h��/���b2�'���~Q8�����_3#ڸZ鎬������v�R����/������!n}y���q���U���Ji8��>|�(�O�*8$��N�S�)37J*uc�A�L'{Z�˗D�6���l ^�V]��}R�wX�Ղ����|���P;H����!n}y���q���U��C�k�j{�C�-VB�T_3#ڸZ鎬����/���B։!��a�i\��[����<��z��}�Q2�+�Y�%⤺���b܉���i�kL�5N�6�vg;Je'���Xw.9�	3�/���jbPhrK�@<,у7G#+��Q2�+�Y�y�J�#z����ͩ^��8k>6s����]�!��	Ǹ�y85�������&H�[&-n�g��U-�e��A�uި��y��Kᷪl?
�A���~[9��:@IE�U��@�ڗe'T���+«7SŞ�Ӣ��WT�j
�I��w��,c�A�L')��7����0�7��65�&H�[&-n�g��U-�e�4o��0����`�3�E�����7G#+�ǟ
��|�6}.�Q�º�F����UD 	mO85}��A�"�b���"v�l��9�4�3J��Rs��@Sf<��orǟD�ui�+��V�-X�G*.s[Ɠ���]{���qi�k��E��z�tP�����ȓ�Z�ܶz��gpӮ�;ۂ��IÙ=�H�^�!�8��-q�@I�2����,��YGQe�.�'n�^0o����y�]���U���eu��<�q{�f��a�:&�>��s~7*� ��RC U�<��y�3�Y�`�'n�^0oza(���D^�=�Q����f̫zjI!JN�K��J<W�f�ӊ[�k碝{l�f|�ό���.�Xu��k ����ͫ��!n}y���q���U�s��Ę�5������:<��z��}�Q2�+�Y�y&��{)֍.�F�_3#ڸZ鎬�������(���n�Ak�����~�s��g��U-�e�4o��0���)�XGG�č�Y���S�)37J*u)T{6T'=l�o �<�����!n}y���q���U��C�k�j{�C�-VB�T_3#ڸZ鎬����	�+9��\��*�J�Ϸ���W<y�׀%\ f�Lu�m�WT�j
�I��w��,)T{6T'	W��^$k�i�kL�5N�6�vg;Je'���Xw�`��	����%n��WT�j
�I��w��,)T{6T'�:���N3!!�[Oj8�6�vg;Je'���Xw�j�7���`]�n�p��owђN�~R�wX��.Ï�� C�(��EZ �:���Q�6�vg;Je'���Xw[�k��x��>�h$G�����=����(�
t��Y�{'%s=ͱu��̦�"�K�b��Ub�ۙD��"X��[�`�L�i�AKd��y c��$� u�r]�D`�6�vg;Je'���Xw�j�7�����G�W�̩c��@PǨ�o*� 7�v�ԯ�`�L�i�h�u��S/Y��P��4��6�vg;Je'���Xw��}�m�kx�-��g�S�WT�j
�I��w��,���|HH9M\��e2��p-!]О,���ۭ(��~T�����DM����p̢M8���2x��Sd[���]�LBt�&� LK�a�]G��wi�bZ��b�Bv�~������]�!��
ך��T�y��9/���`���6j��|E\0�*�W�ӝP�|��].��'���XwN�U�R��7W��!���{l�f|�ό���.�hM��{ �`o����;v�~������]�!��	Ǹ�y85���*�t�<�uծ/�,0=]^	�&������ *����h�(���e����{l�f|�ό���.ӂ����|�*3d��'�|��].��'���Xw�`��	��d^�qT�b㨵�֯��ҋX����@�ڗe'��.�f�8La���R�l�>D��(�
t�ژq���U����Q�S^��c-(���X$�{�b�@IE�U��@�ڗe'AKd��y c��"|�썥��9�dMbZ鎬�������(����l�`�n�>���/7R�%�T�\ �̈́��շ+���eq(1p <�r�\���ҿo�"aI��w��,)T{6T'8��������)��[68k>6s����]�!��	Ǹ�y85�Q��%s�@�zl���y���/7R�%�T�\ ��&M6^�Jm!�<��6�בa��@IE�U��@�ڗe'AKd��y c��$� u�r]�D`�6�vg;Je'���Xw�j�7�����G�W�̩c��@PǨ�o*� 7�v�ԯ�P���<e<>\��p}�	��D܂�A��W8ƭ�I�p\�WBQ�,LA�lή[*%��J{�+�M�( �����+�@{fT�1�߽K}��׍����}0�st&���\�vūx`��:�,�qo�,ܛ�	��|��	(���zL͊�q���19TH��@���U@���:��F���V!���IÙ=�H�i�͒/e���@	Q�č�Y�����&��J��7l�����x]X��I��S&ϊ�fݘ���GaY�����'�u���vb���@���8y�)��j7T$�S��^y�8�>W��M:��2��mc[�o�v�~������]�!��%��rSe�uF��θ�l��o��H"
�ҋX������S8�/ #O�)�t_-Z��T�\ ��
]�T��i}3�J��J�*��:�ҋX������S8�/ #O�)�t_-Z��T�\ ����)5!t�����rl���בa��@IE�U��w�B[��lQ�$�k\_x���� �Kl߯l�A�߹z/�=�I=���ۉԮH���v^�n���!2�ͨ^��e�]�\f��F�K͕[y�������o��C!T*�q���U��s���+M���9$���]�!��:=�1:��{oAS�i�<��z��}�Q2�+�YɁe��b�ޥ�o��C!T*�q���U���X��u�����
L'���Xwݩw�_���
���)�b���"v�rJ�IaF�<��T���:�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��Y7�u)S��r)�o�$C��c��(r���2r,~�oHZ��S�b=��%'�_��z�������ZI���~���U�z	��ߓ]�>k+;��5�k��y׽)N�[SV��˵��W�[4�	�}���^e@��V�i�I��Mֱ�H���� 5+� ��G�|��8��\n$̱̉���ߊ�,�'��.	&'Q����^�[��$*�¹�>D�� ��;����=IEw� e8�~�����0�H��OR�JO��V�RDFR7�h�Qf�����m���t���S�����ۄ؈��k�;4 e8�~���zR���bp;EK�6(��Mށtd؈��k�;4 e8�~���zR���b�W� D���>X[V��kC��8��h�Qf�����m��u&^3X���W��'LC��8����9&���"E&��� �����祎〕p�.��G�+-�q�,a��Z�q�,|�)�֢-du��~
�^^���X���v'�!��	�'�L��OR�JO����9x_�+���{�����w)�0�7��65�'�2%q{�f��a�eSܥOH�?�o>�q-7�� ��͌4s+�nyo�)��9��>x��F�\��Ɲ&���e�I\f"�	-7���J��ڮb�'���ߌ[R)Ms	[��c<+0.��Cҷ��eZ���hP*�g,�5�TzJV��šoLw8:Q�{4�5�Y�w���Q�`�B���B��!_O��Usj1n�1a�m�O��]�lEGV`2�s�f�6��5:xt�mdy�-��g���?�om��;���B3t�yL{�2{�=��E�Ծ�V���D/C�H��a�}8n�dY92"�f1�p,`V q��~�'�<�y8|�g�֐�o30�@Cq�,|�)�֑���w1�'f�wR�l�U�X��Ŏ.�/*��9J�]Sh�=�}�2����X+#��;ϫ�7�l�h�Iv01q�k\ ��e١g.�ե���.�U� ]��ɦ���2'\�d�����ca[�2&�;ϫ�7�l�h�I]����ljrk�� aD$O�x�Q�Q�?uG�Qy������(=2�u��s$y�刢0�]���,mxX=��uZ��הX{\�IV!"�:���l����R;5B5Y+�N�#�ɉ� e8�~��;�r"��[e�A`�M��V.�g�.�ا�v���}�{��<���#:B�Oy�~�R�&�����h�Qf�㷝�u!����7��=�B�z�\޳->��DV�RDFR7���X�A$(gKk��b�~)����n-Yg�yi��v�{�a�,.��/l8,�H����I��'��$�R�n����͛��W�c�'n�^0o��0I��I��'��$�R�n*d�c��n�b�a�JHn��z��`�B�92Y��^@!�PsgD@LM#��aPSp¦�5����`KW+X�~{�\���M�
`�t�啷�q{�f��a�I�4T�E��EMU�YG;] ,����a�� kF��4�	�}���^e@��VQi ��M�r��VYW\�z��j4��Rm�Ƈ��ݱk4# ��}��6���'n�^0o��3`r{�@~��6�% ���+a�G3�u]��;�LaP�'���ߌ[R)Ms	[����a�k���� v�D��qz�L<�������r���aM"��N�߄�4�X�)Х��Y[�P��)��\�v��N��V^���VB��z_��q�s-�#���[�"yd��N�}�g,�5�TzS�@/{�&ӧ�&��������s�����	)��59�M$#�fJ��<���6ɺN���ߙ߶h��M�k͝���:2�_]�5����`K�A���Q������;e5V�]C���[���?S�*���X:�*��ܟ���Gm_n��!$x�C˭oϨ�{�ś>���0�qU]�Z��L<�������r���aM"��N�߄�4�X�)Х��En:ъ�7k�%����x�ݠ�oY�1�O�vf���Wi����y�:�~%��;@6C�leKWa;.]�n{l5�z�}���XH���E>��V�Q4�:�^���A~��j.o�c�\.U1+]���H����XP���,#�N�MĐ�r�
���k�û&�l0�3p,����Ѓd��g,�5�TzS�@/{�& S�t����� �C��b���:� ߬����c��1���8}�Ͼ'���ߌ[R)Ms	[��l^V���
���*
�I��'�yۨ��~���CǍԽB�Z鎬�������(��＂��@ê�]���P�.�a(􆿳�tP"7��%�j)���������I��'��$�R�nL��C��&k-���h�����Hb�zL͊�q���es�1U)���\+N��&�L4⭦�����.��r�3�������r���aM"�������4�fN.�����?ׄ/�L	ACDCx��-��߂��g�K�
��$�~ȣ���XP���i�7��BQ���b�ǳ�LU�C��z��-p�Jj}Ѯ��.�x��W+X�~{�F(�E��p��+ᕮ��֫��XAьb2up,1�-�Y�}�ƈ�L�i����uZWC�O@�����K�Q����
�?<J�!�Ӑ�O���?�]�!���1����mB�8r\V��P?��������]�ٻ�q���U�pzl��a�V�RDFR7��/
����X?�WGc"�Ee�6;�ﻋ-���C�M��N�����ıψ6P�p�HZ5X�vZ��B��=Y��_�n������K�Q����
�?<2�,)�<xE;KC\�d�٣��c�A�L'M�Kc�I؆h��l7^*(��oD���g��U-�e�۴WLFo����|ՄT�٥��T�A��ˮ���nrm؊(��~����p�d~c�s�����_���&Y��V�c�	��}��/刲�ZT�p�n�ͩ���Z��]�!��	Ǹ�y85�L��0�͂=��«hj��I��Ba(􆿳�P��AK��hx��W̗���%��Aс�^�r2&����Z��beNY��;�W f�Lu�m�?�&͜�ﻋ-�����S8�r�:-�����`y����{�-�;���0�b��b2B`Tz�����mj�pzl��a����G�/�Sx�lޞ�ό���.�	[ZZ��g$������B���؈��k�;4��K�Q\���q����� }v����5�ź��=Y��_Q2�+�Yɂ�rS��9�<T�4�B�8r\V���6<p�W�\��I���Z鎬�������(��＂��@ê��uծ/��T�\ �ͺQt�v�����bC��nrm؊(�pzl��a����L�Y&Nkj�w����X��'���Xwd�n]N��l�`�n�>p��HM�e��`y���k�)T.^_��ˁD�wE
]3b�J5�e`��9�'�E�Jg�ˏ8[$0����X��'���Xwa'�<� \aXԳ�>����
�?<���+Ɍ�pZ鎬����>�ȬGX"RB�8r\V�7��G�����a��@�_!���?GQ�.�!��kw2k����W]�Xscr�2u�蜍6�����=Y��_<ͧ�:|x;u����f`�	#���/HG9�G�O�}?�P|�z��������>u~9T���l�FWv7��ٌ���eT�]�!��	Ǹ�y85��d!+��T�"���N��MY�5����;�
�(NJ0�������5�e`��9\�RӲ�I�j�?x��$�*�фr1���F"-�`��8�4͇��U�tJ������8`N3�r%C�c�zȮ�P��fhH�{u��w1j��a]��R���YC�X|��K�Q�B �n�6ӌ�Iۏ��D����1l:>�<��ﻋ-�����S8�bM� 2)G��8���/�.R��O�vb�
5�[�*ؐӘ�� ���2��K�Q�B �n�6ӌ�Iۏ?�WGc"�Ee�6;�ﻋ-����2�77�EV�RDFR7�|u&��*����is�'ח�B��&ʧ��Qe�*u'���Q�@��߿���A�U�u�;�����K��[��f7A��(�n����%HlܡZ�0~���/��H�)�`p�ʘ���>����0ʉ�}���Nu�U|^Cf%���>u~rۤG�#r���#�g���#� ��>�%�*/@D���uL�-������������,Q�o�Z�Y�z�r��[��7���9����_X3�G6t�T>�"x��@׋8FZ�±��m���*�N`v��W#�����^5J_�>Y�{'%s�6F���y�g��U-�e&��B�v(�T�nf(\5fٜ#�d���4L"�#�4p`��k͝��5w"^	��)׺�������Jhפk������d�٣��Y0����k׌"S�0Q���g��M7�mpU��C����$j�@�����x'T��p��`f6	�FWJ�)T!��=e�����1p�u�]�!��mi��d/���l�؊9�p'qc�	��)�-���a�q���l�pzl��a��yu>ý���9,3�<�P 3�'���Xwwd�t�"��*蓱Wxi��U}t;#60vn1|3�!������y@���ıψ�|���!��M;�E��C��'���Xwd�n]N�z_��q�s-�#���[�3��z�/��^�V]��}R�wX����K�Q�	y��J����9x��iҋ������	?�4�]�!��	Ǹ�y85��NÍ@�xx�rDc�O��Юlb�'r�����8���/�a'�<� \�/刲�Zh�X�/�.B��p�	Z鎬�������(����ｗ��u��?��Q�&{��8�aЦ��W��Z�8���/�a'�<� \aXԳ�>����
�?<ТKH�{?PkF{����rs�i��=29��aDRŔ�rUq��ɤa��)gΔc�ȷB���������ȓ�iӚ/��MN����!I/�������A��X�@�5��6�l��s�����[� y�~��ż3���F����T�O�H'�J�����=<�HI����>�W�_=��0���̏�u�=Cm�v4��61��7a	�����Y�
ɸ�oƴd��t�'��9ܛ�	���V[�+
�l掝�K\m��U}�	|^�׽R�s�DH}�_z�9�E�\����8�i�`!31u��Dfd�W�ϛ9����ɧ���7�)a���%}D�����!��g�-��\��OA�=�~�]��d�Y��o�6�֟�Zl��a>���(�WI�;�_�	�t쩖NUD60L����L�Y&#t����n�~����p��l�n�Zl��Ͳ�8�3���!��@HW7��ո\����8�L���9���D�K�X�Re�d���L$�ѸT���C6���$73���'���)w�i����0\p c
N1�V&�����O�qTkή�Ádo�dvAg~�r{m��<�te˩���.|��f�ͣŗ�:���+"�9���B�I:׷�F!���H�v�!���y �谝��X�e�F����To?��m\Ӓ�qܛ�	����%��1����ї4�z��pU6�M�S��2�{��΂`g�O�.UT��"[�(V�0r�����K�9y^6gVW���%@�~� ���I�����+����>�G0n�>���@��3y
�*����zEK#�E��Ǵk�?H�$�IX[��O2<������ #M�)��u��`�|�&�#�E�d��������y��Ld_���1[���K��&�|�G�2I�wp(��C�712��}ǞK=<^��`Y�F�����I��#��
Mcu�T�M�ڤ [�f!�)�X�j(�� ����n�
_��q���<�{�!���"�ֱ��R8v��j.Z��$�sӢ�]3�����c��(r$����Gd"��U"�̩��k&Q��8�'��j^ҩ#��u1�L,Jz�փ�G�#�j���Օ��܄��� MF�����N6�@P�q�܄��� M<���Hn
V~$�A��w;�Q�40N�J�O��~�Zc�ӭ��Y)�/����7r�Tة��n
V~$����6��O��=?u�gt�DY��b�fc$��bӴ�"�6j��8rW��N�Lq���Bl$P�ĝ����v�pmw�97J�L����߾�'w��I�MK$YҦ���Sӈ^t�lHn.�����:�'�׏�����Mx(�i��/R�������a�U�ے
9�GKP�2�����Vc2�����Vc�cRq>h�,���Ξ�I��CK�8�:R?+��7� 9�GKP�2�����Vc2�����Vc�cRq>hLV�4�ұ��ݣW�](������(���4,e�b�����E(��6���s�
>{J�s���v�1���W�-wP0���wdo�6�����Yw��-�a���v��^�o�A�r-�lu���D��ܒmQ3��TO�$=�Z��ͯB��ooF�!ݒ���|k�g���鞨��k��/����h#����f���7l�"b��"@��}Q�V�I�o#��� �߳G!74/����:���N3!��u������[�)"��H��2���r���2�lW'+�Q\9f��qb�Naْl��]�Bc�jv�Тkmt����]$�﹈�i=p�f�[��iO\
$�*�_���C_�!/XW�������f�w`�Ӫg[���+>g�m>�`^���t��˳���f̫zjI!JN��=ީa)�!��ZB��,�Ӏ(��[��B�IxoҢbu�ߞ�(ɡ�>�(}%@��7�����3�!`�mL�b�-G����� 5#�3j��dǑ؆�!��ZBV�RDFR7��/
����X?�WGc"�Ee�6;W�S/f��e�WDv�b��h�Ӆ��x��-�"E�3�!`�mL�b�-G��'"�}�u�>f��+����ȗ,pr�B�,{�6P�p�HZ�$����_UX����;�eL�(j9W~�O�N�H��!Kp|��+�Y�G9�$�#o�]�lEGV`2�~8ถ�#�T�!�K����l�?),���'^^�ȴu]���ϋ[R�S�/d]��iTN�m6
�DR���^�h5���G�?v�������6�`�۲r(ϗ���	X!�w�H���-!����
9�B�ݔ�]<�7~�����M���0t9X�8�ޑe�ռ��@�[OJ�k��A�,����	�|ϋ[R�B6Ji���5t��vRTɷ,iS���tk�A�,�4���/,��YHiJU�m6
�DR��shܾ }���R=6�&���\mИ|��,���xoqUioέ����go�+������t^���\�}����
�?<l
b���p)�i/j�ooF�!ݒz�]��b��R�[��ݚ|]�dT�'��7p:��g��U-�e�$�R�n����͛�v�!;��w��ٞ��/>x��F�\��Ɲ&�n�Ak���
h�q}lx"�fu��ė�P�"Y��^@!�PsgD@LM#��	7>��5t��v��M;�E�p)�i/j�ooF�!ݒz�]��b�p�(���J��� �C��b���:�벩��Y�W+X�~{�\���M�
&��`1�d!j�e{�~��j.o�ѱ}����SǴ�`"��x8
X	:J�/����CM��ߪ���W0TZ�>:��aB�e��m�|�+��?�d���&����;�Ӏ�S�/�TX訬ȫ�A��R=6�3W[��l��Ȑ�Ӻ��L�~�y�ю�?��Q���FQCs">*���։�s/�~��ꔖ���q�b�-G��'"�}�>�*�L�ʽq��4ȇc9 r�e�zf��7~g�[�!U���5��&<��iD�H	�����
�?<�09%?�3�1tm�/Y6P�p�HZ�/?�?6ר�`'֊�D0r➜~yٹ!5�j�B=?��FCC3Se�� ���� �C��|$T��!��/8^b��w;��|B���?#�+~���V$��]���e��=���)D�3����hF���O}�Sa1����D�3����h5x�<*�f�R?�6��'�|,kW�A��ˮ��V�rsSRą�3E���q�kGQ��l�4��H���EO�{���V����SC/���d}��[�ƭMj��-2/��2�����Vc2�����Vc2�����Vc2�����Vc�C0�M��VL��*5�tK�h�+�lX҉~k�X���2�����Vc2�����Vc2�����Vc�cRq>h�e�B��m2��+h�ˆl��=�j� f�Lu�m��)�u������k	D[b  �H�,3�V���C��4c1�~v_��s�֙K��J}L���E��1��8f�؇��*-|d{�A��>���K
��c-(��z@�o	�Au�_�\�Zr�m��n��&�7a	��������W5�\tCՌV�����,����_,�qo�,ܛ�	��������'�3�$ �#^�Vn���v_�"c�PƐt
׫�J��!��l��[�?2^�9�ԋGw�����N-6�m~G��;ؔ�Z�	���$�R�n�6Knr��X��-�`V-u9�`�T�}��K��b�!cIh�{V/�_��د��� r�	�����ވ�'��Ǵ�X�)Х��㵾�Fz5��F�g,�5�TzS�@/{�&qóf�ǡ-�#���[�"yd��N�}�g,�5�TzS�@/{�&�_��ƊH~��j.o��)����n��3;�í��>x��F�\��Ɲ&�O���EWI��X�)Х��B�O�n������r���aM"��N�߄�4�X�)Х��=�\2�lFb7�v�ԯ֗Q"t��������20�3p,��x��δ�OUioέ����vЧ���ܔ���1������f̫zjI!JN�ߩJ�9�h���X �Z�^6.���6�����X�V�RDFR7��D�
p���kg>�[OH3=-��7����@�}z죹`Zf�Q�@��߿���A�U������W3@���ӹ܄��� Mh���X �����R]Y䅀]��uxe!0�K�r����h�ᮛ�ڥ��!���α�%�����,����۰5t��v�Â�&�V���do���;���GU)2����x�w�Xb<������
�?<f ;+/���a�{��t�N}�}���
8	*�?�*1�#�;����הw�u��Lj�eS1����	jp.�����w�r�^���1n���6�|�+��?�d���&�<��Lio|����&���o>�z����
�?< *\p�+�����&�䐛>F�%<��7X�y���C��"�v�Gf�4�ͻs�	Õ�)X�J�go�+��Ŵ#����#g�k��5د��������z� ��!���\�_�Hw޴]�HB�Ǉ�h FS���Q;�im���M:��2���ӳ�Y�
��e�W+X�~{���~�G!U$Y���-X�G*.s�FÖ<^������V1鴥�`B�g�c0���]�.�Аv�മ#F&�8�k�<��~wD[����B<:���-65�H]k�'���ߌ[����65��F�g,�5�Tz�o b�ўw�� ա>x��F�\�=�5j�˛ݧG �ŴP��Cn**�8����>x��F�\��R�>�v,0=]^	�&bMydjpCb���z��>x��F�\.��0�3�^�XKS�*���X:�*��ܟDY~��;e5V�]C���[���?S�*���X:�*��ܟ�M����یӺ��L����~�pP�R���+a�G3�u]vj�[4BǊ[
�}3��C�X��z�f��&@�ES��Hس�����L��S-������%E�X]on�ǚ�e�|��ooF�!ݒ�N�PP�}hU��xz�J|T���2�rۤG�#r�X{�"|Ӎ��5����'�)n�J��ָkd�vu�Z��F���˺�Q���|�A��^W+�zN����!��ZB��M��7X���@l�<�){:��K�}i� f�Lu�m���Ț����WDv�b��
<wͭu�H3=-��7��B�>�93�!`�mLy��[�b6W�����E,E���Qk!��p�1C��'�mw ���NoǢ R�*�߾�'w��n�Ak����h]f��Q�4���܂>\��p}�V��	��yv�ʯʗ\:��{�ϥ#���,�+ f�Lu�mo{�K۬��%�^O�����k����*�A����tz-�u�O2"k�C��C��v�Gf��$�R�n�m.�>"���F?Ur,�;��|BD�s~��'�B~�Ǎ��d\F��.��#��b�]J2�d1Z� f�Lu�md0
\,FQ0/zﴚ�F��Mu��M@�1���ۉ�8j1��ْl��]�Bc�jv�Тk1�%n�@��V�����<o�nïi��PL{�ϰ>D�c�lQ�(��Q|3��'�3�$ �#^�Vn�����'MRmHX���y�XZ@po�ͫ��;���^hq��:�V��ÑR ����*��Y~��`�J�(��Q|3���ӳ�Y�
��e���`=����wJ�G�����t �/���7R�L��_���	��f�!"����}�Ay0Hb�Z'�2%��5��v�o4�	�}���^e@��V�v�AZ���F���9�@Zd��`�H�&���1DV�H��~ж� ��%lsσw�kz��ՁO�#dh���X �@B��ї�ˏ8[$0��ґ�po*��p��U�d�K��@e�|�\����t	Ma��S��W�l�l���XU(�a� '����X�*N/�p��m�QKӲ�g����[��밼�ۂ3O��R-S6�o8:4ڛ����R]Y�bF�B��/�
k���6<p�W��08&o BVf����aUŪ|u�?b�L���dL7A�k�6���rx���g����[�=�.��c�Z�&�Za
�	?F������������76�܄��� M<���Hn
V~$̀w0��b�#��6/��������\n0�8�_+ӌTkel$P�ĝ���Pع����ɷ_F�!���Fi����o<���H@w���H��j�Ï��	p8,3s"�1< y��Xscr�2u3�J~��k����VPYUt�\����Sӈ^*1�#�;�e�*[�9�������;Ϡ������`:,���"�&Es�];i��I�x(�i��/R�*�W�Ǹ!2�͞nOY��m����e?�d���&�V�RDFR7��,�p�HO�]N�&EЏ`��S�����@*���k����*�A����tz-Ղ���g�����ܱ��KOyTg��q)W+X�~{�ւ���z�D�JM2�_��s�֙���^K��Xscr�2u0�DWB�=�<�^����,�ǰP���Mt&d\F��.�����
�?<f���BG�ܕD1`D�Z'� �Y�2�����Vc2�����Vc2�����Vc2�����Vcl��w&� AJb�!����l\�:�D��82�����Vc��g: k��2�����Vc2�����Vc2�����Vc2�����Vc����1s�g�qL7�[���V�1�RR�,�*Ǚ62�'���v�����̣��4�#g�k���ح(��? "a��N���AI1���Ѷ�0�rۤG�#r�X{�"|Ӎ��5���l�1C��(�V�RDFR7�t�+37/���@��.ڜ���,�ǰ6y����m��j��/]/�֍r�
S7U��ކ<&�|�����l1� C�z_��q�s-�#���[�t
ZZK�z�f��_��s�֙���^K�����������f��M���\��E��U���}h��R�Q��=f׿�������!N�2��_:��y$[|�h���X ���������R�@Q��oL젡�q�FƈxN��b�@����F���9�@Zd��`�H�A���P?�Ӧ��Z��z=���� ��i
E��l�1�ԀU�܄��� MoE��cFl�㬲C^e�|��ooF�!ݒ�N�PP���Q*J�<I��%����b�md��/����h#�`z����0Dk��v�A}-������Sb���!��ZBu��w1j�C;=B>���h��śa0��#���N��;�Ż���fx�ZT���2�rۤG�#r�X{�"|ӍLQ��}S�r
�w�f0{��
���S���B �n�6ӌ�Iۏ�xA�)�X�QP3 R � �9D^��kGQ��l�4��H���0�0�h��#g�k�������h=�I����KI�R�'\�RӲ�I�j�?x��0���x���
k�jh�Ģ\�RӲ�I�j�?x��0���x���Ϛ�c������锴�;��|B`���m�Q�@��߿@
9�"/�@��Flp��u	����� �Q�c�C;=B>���h��śH���_�/Gq� ���	z�Z<��zUD�3����hY���v`?�d���&�W�!�
��i�!�� .���AOXu��w1j�C;=B>���h��ś͙��V�����O��Q�@��߿@
9�"/����+�,M�A����2��O�c����X�)Х��1��1�_[���Rm�Ƈ��ݱk4# QO�jv�k���锴�;��|B`���m�Q�@��߿@
9�"/�}�Cr`�r�u�fv��c����)�f}Q���h��Cp��I����ۂF?[B*��B �n�����7LH�D���Lxx�rDcѴ��B�66�� �r;����9:�B��B�
/Sq�\�RӲ�I�j�?x��0���x���F�s����H���MO�/WOF;�Z宨¶J1�j�$�R�nL��C��&k-���h����k�S���S��+���Ã8�4��Q>�u��w1j�C;=B>���a��$���}�����j�s��1B"�A�`�=�ȭ^0E���^��0�$�ð��T���^���Y9T���l�FWv7�WIR�Q�a�vU�D�}�FZ�±��m�^p+�b��>CZ��p]�/HT�Y�[V��M*W+X�~{������Ll.�v.���ƶ�~b�!jS&�7G��~�޷Ζ� �1�f����y��$*T`�̍"�����{����r�&�O��p��D"����#CK���L����E`���rw�&�z<a��N� φ��<�6����s>'FZ�±��mJ^k��ô��Njr�Ú��9�2�L�B �n�6ӌ�Iۏ?�WGc0���x���"�Ee�6;Ps_*�GqW�w��fD�B �n�	��c�n� �Q�c�gt�,�$����;����~Ϟ3-��U�C��z����7��j�5 �X�T��8G�<e/v���x?ߕ���Z�רXH�b�:�&�e���F30��	>A��jӁp=o0";��@I�ȅY�I��;e5V�]C��m͡r��b  �H�,!ԱX�|�4�`a���O[H5�NUAV�?���qR� ���I�S�S��|V�ؔ?%b*� ��~�8N|��7�'�L���E f�Lu�mf׿����q�>�Y�V�W|�B�I:׷�F׫�J��l� �[��׍��������֡�\�<7�X�e����]��m�n������"���P�`m��';��?2^�9<o�nïi��n�5�F�^hq��:p.}Tp׸I�H/�v�6���l �{�!�e���,��`/[�f;q�s�|54�
1�RR�,�*Ǚ62�$�؁�۟D�$0-����G���y^Iiϫ�Rm�Ƈ��ݱk4# �W�ڋ�{�K�b��z���Q$�@�xx�rDc�5��ja~��j.o�c�\.U1+]���K7v�14�~�Xo��X�Ü3�^�XKS�*���X�#Gw6��>�u���g,�5�TzS�@/{�&>ٮ����l����B}�S�*���X:�*��ܟS^01D�F��l�ꐘq?U�C��z����Ջ�/Cp�14�~�Xo��0���8Ô��A��xq%�܌Ӻ��L����~�pP�R���+a�G3�u]V�`���.�;1?�[F�sp֟kh����aA�h�Ӆ��x��_���wg�W���'h�]^9����]I�r�B�,{�6P�p�HZG"{�e
Y�;���GU���|k��v·��\�RӲ�I�j�?x��n���Ϩ��`��X~���t���s��Ę�}��U���)���w^J�b�=�P�K��J<W�f�ӊ[�k�T�"2o��3��	�3ַheJ��D��v·��\�RӲ�I�j�?x���Ț����WDv�b��
<wͭu�H3=-��7��B�>�9}�����ņ�a�t��S����k��l#QF�ky��.�"����
�?<�U
��ڌHs�3�:����k=5�Bmy;;���0��0��}�<��WX��Yб�鮔C��c����U��\JD�@���:�ox㲐�a�A��ٞW^�TG@|3sИ�c�2Xy�WwꕶI�j�?x���V��&|6��7|�#�I�ȅY�I��;e5V�]C��m͡r��b  �H�,!ԱX�|�4�`a����!�T�.�xkx U�_@�Ǒ�\�J;&�w��9�0��0��}�#���,�+v"���'���mN��"M�S�Q;�im��ɝ\�!2A�X��-�`V-u9�`�$�E\�<xx�rDc�O��ЮlbՐt^UYܓ$�R�n�9j�ʛ��!"����}�ܡDi9#_� 4j)$�|54�
1�RR�,�*Ǚ62�y��{W(3���P�5��$�/sNc]N	��14�~�Xo��X�Ü3�^�XKS�*���X�#Gw6��>���s�Tѡze�áS�*���X:�*��ܟ�jJ����d_��=
R��Ǔž'���ߌ[R)Ms	[���$š���L<�������r���aM"��N�߄�4�X�)Х���އ�)U�� 6F�GXI.����Gވ�'��Ǵ�X�)Х��㵾�Fz�������p����c��1���8}�Ͼ'���ߌ[R)Ms	[����.k+#�Ye�@[o�����20�3p,��x��δ�OUioέ����vЧ�����~�;����v�������d��`�H�窝�0k�����h4c�=���� ����%E�X]on�ǚ�e�|��ooF�!ݒ�N�PP�����%E� ���1\U� ��Z�!3Bmy;;���0��0��}��yǯϷm�{Ξ�\�s�a�{��t�x�X�ڹ:}��U���)���w^J�b�=�P�zc՝RqV�H��~ж� ��%lsσw�kz��awf��!��ZBu��w1j�C;=B>�)3����Հu���%��K/�(R�����%E�"�Ee�6;��v·��\�RӲ�I�j�?x��n���Ϩ����t����E8��5�:{�#�	�����1p�Z̘�Rs8�P}�����ņ�a�t��|��[}��t�G�h�J�P��g�V��	��y���rk���&�e���F30��	>�`Ldk���hi���D�;E����� p����勃��;FZ�±��m�5�9�59���#KB� ��~���4M̍����Q6vmI/5(Q�g�+%f���at�)��d��X��WG ��օP0��p���Z۳
0.�
rQa���d��{S�u��w1j�C;=B>�v�{���	/�M��7O��4'��7�OT�,�$�R�nL��C��&k-���h����k�S�o���wu6��C�#/�����r�&�O��p��sW��/�����ņ��Z۳
0.�
rQa��Vf!�q�#k�˟ܒ���靤�}OJ�1���۪	�}a4�����d�I}��Bmy;;���0��0��}��`��X~��c��/�^N��P�vJ}���j�s �O�,R?����>̞f�2-��������)�>�#��FPs_*�GqW�w��fD�B �n��Ǒ�\�J��0aW��/�:�Ȍq[�=z̲��\Tb�:�y<H�D���Lxx�rDcѴ��B�66�t��3>L��Q���_��s�֙�ɋn�ŕ� �U1!e��`����A��jӁp=o0";��@I�ȅY�I��;e5V�]C��m͡r��b  �H�,!ԱX�|�4�`a���O[H5�Nxkx U�_@rJ�IaF�<�����J��
lR�1_��-�/<����ж�Z��9<�)�$��@�e�3e�����orǟD�uiM���	�f��DriU?�7a	��������W5�\tCՌV�����,����_��*���3m��U}�	�2�G�Ml\P�O����X�e�.ċ2o�0ad&(C�#�7#^�Vn��@�P��.�/'��"���P��_�}4U�&�L4⭦}��-�ӛ�!����X��-�`V-u9�`�$�E\�<xx�rDc�O��ЮlbՐt^UY�l�;�w���h���X �2�%͝m"�14�~�Xo��0���{K�e�٦�A���Q������;e5V�]C���[���?S�*���X:�*��ܟp`��2L��14�~�Xo��X�Ü3�^�XKS�*���X�#Gw6��>�u���g,�5�TzS�@/{�&>ٮ����l����B}�S�*���X:�*��ܟS^01D�F��l�ꐘq?U�C��z����Ջ�/Cp�14�~�Xo��0���8Ô��Akx1���CUioέ���K�IE�����s����i|StߛE�������l��;�4~���;A�/'q��������|AW��0���������L��S-��N��3S��%�j׾���~�ch�B�_�+�)���&���/N��3S��%���|k��v·��\�RӲ�I�j�?x��n���Ϩ��`��X~���t����z�+��p�,�#�w{:IxoҢbu�ߞ�(ɡ�5b��-����|���kJ��K�}i�e]y]�g��!���α�%���ޣ�`Zf�Q�@��߿Ur�g�g?�E��6�)�b��N��3S��%)2����x�w�Xb<���B �n�6ӌ�Iۏ?�WGc"�Ee�6;3��+�W�Qk!��p�1C��'�mw ���No��`Zf�Q�@��߿+��F�+ƓƓ+�>\'��%9j�m1�H���W�w��fDrJ�IaF�<�����J��
lR�1_���KR�h�u��S/>��ᓺ���)���IJ��%���R~�hRU>�����r���aM"��^��J�Y�y��{W(3���PYV��
��;��|B��w�>�b�����(6ӌ�Iۏ�=]92Q���B�װEl��9�4�~�ۉ�w;��x�l��1i�t�U��D5l�_�G��G2ŝ,\�=U�C��z����1��t!U$Y���7γҬ�,;r�mR-AFe�oU�Hh���{|���?�}�h���X �ݧG �ŴP��Cn^�\���ĉq�p�F><1���*-�RԚfވ�'��Ǵϴ`�-2c��ҭ��'���ߌ[��83�$^�<ĘX.�
R��Ǔž'���ߌ[R)Ms	[����80���Z%ӗSu��z��j4��Rm�Ƈ��ݱk4# �
)�������4�a@�B%���O-�#���[�"yd��N�}�g,�5�TzS�@/{�&�<�?�aޑ�74i⯶��r�p@iV�g,�5�TzS�@/{�&rM$q�̅�	5�8aw�1�RR�,�*Ǚ62嫫�Rm�Ƈ��ݱk4# ���M3�=F�8�&��A6�k�#��.���t�:�6[��j;v��0�3p,���#ip��(f���˶HyNL���&@�Ex����MԲ���d��#�֢W�p�
ͭ��]I�r�B�,{�6P�p�HZG"{�e
Y�W�p�
����އ��&�nP{�B �n�6ӌ�Iۏ?�WGc0���x���"�Ee�6;��|fa��^4/��?E�l�1�ԀU�܄��� Mi�@�ZZle!0�K�r����h�ᮛ�ڥk:j%]a6��w%e�}�����ņ�a�t��T�b^ �%K!�Gr<�*���do��W�p�
͚�� Y�b�4!m4�UVu��w1j�C;=B>�y��[�b6W�����E��t�6��B�O�
B��$��~a$�B0�C�Z���}�����ņ�a�t����>^��m�b�����(|oc�݇2�۪	�}a?�d���&�����[1o�>��ᓺ���)���IdiVbL� �?�&li\�]�(f�ݗ�oFIcfxah���(f���5�r*Iީ�V��F�-���E.ƠGCe]y]�g1K����4�0 L?�b�=�PXu��k ��Н" )\�RӲ�I�j�?x��!��=e������9?��k�f��a3/���%-��`Zf�Q�@��߿+��F�+ƓƓ+�>\Z2/ڇ��B@�L�q}�����ņ�a�t��|��[}��t�G�h�J��X�����V���+���Ã8�4��Q>�u��w1j�C;=B>�v�{����o�kQ�@��g�0�u\=�~ o8�1�R�*���M�,������3~I/��\]=��"�ԭH���MO�/WOF;�Z宨¶J1�j"�A��"�Bmy;;���0��0��}�<��WX��Yl�3@\h��`,9�H�WF�)Urx�$����5B%���O�����4��_���e3,��V�.o)�B �nʃ��#�a,n�cqgF&tS�D�H���MO�/WOF;�Z宨¶J1�jn�ţ�Gi��(�V�ܼ������A �׏�����MFi��|��wØ��|���؀.ņ�a�t���EF�w*,�AMX��Qm�"�����{����r�&�O��p��	>;�́�^	�+|~�tݧG �Ŵl�;�w����X�:�{������,�ǰ6y����m\du��Ԙф�g�`#����1s��
��TH�����ℇ[���V�1�RR�,�*Ǚ62�'���v���Ɉ����zJ����O�.�#g�k��S��OP�hE�̂�(}�w��u ��8E�̂�(}��[
�}3��*���1���&	��
!�N<�%JW22ᮛ�ڥ�m��k�p�U젩`#ߞ�(ɡ���|E\0�k+�xj�i�S�Eͩ_[Z�g|��ՂU��w�����yu>ý���9,358�5����Н" )\�RӲ�I�j�?x��$�*�фXrt�&�m�����\�~FZ�±��m���*�N`v-��DW���vU�D�}�FZ�±��m�5�9�5��$*I|���؀.ņ�a�t��S����k��l#QF�KI�R�'\�RӲ�I�j�?x��n���Ϩ��`��X~t����_K�@[�_zβrrZ�0m�\��k^��=7�-�u���iq�*C���z�ӛłMjή[*%��J�~��"��ݧG �ŴP��CnM:_A��kg@�"�_���'�>�g;��|B�w����2��G�����#�,$��8�Q�|���!$�N�1z@�o	�Au�_�\�Zr�m��n��&�7a	��������W5�\tCՌV�����,����_,�qo�,ܛ�	��������'�3�$ �#^�Vn���v_�"c�PƐt
׫�J��!��l��[�?2^�9,����_�X��-�`V-u9�`�$�E\�<xx�rDc�O��ЮlbW�F��>���
��Gsp֟kh��/ E�~ (�&��~�~ж� ��%lsσw�kz��ՁO�#d�Ĥ��ࣹ`Zf�Q�@��߿{2���Z�S�����r���aM"����:F�X?�g��U-�e��l� h�Ԉ\&A(`#1/:��!��]ڇζJ������w�����K�Ǒi}3�J���������8?6��תT���2�rۤG�#r,�-�_���c�@�l���=��s�l*O����v=��`x��i��`H3=-��7��y�4K�?���>�lIorǟD�ui9�f?Y�O�`�MϦ��pCeu��|̾?��CG�����r���aM"��h�{V//U���!-�iP��G��\OL^��>%�Нo@���;1?�[F�9��G:([9��qUB������Wi�g���h���R���ɢ���ڠ�Q;�m��j"^�����ϖ [@wPcIn-Hzn�!��ZBV�RDFR7��D�
p���kg>�[OF�ѿa@����v·��\�RӲ�I�j�?x��n���Ϩ��`��X~���t����G=X��i��?Z4Z�7�ɋ������h4c���*R�w׬�H��ŲNGl�R6�.�iGJ�����R��l����FZ�±��mJ^k��ô��Njr�Ú��t���s�3�&$+���Ã8�4��Q>�u��w1j�C;=B>�v�{����o�kQ�@��g�0�u\=�~ o8�1�R�*���M�,������3~I/��\]=��"�ԭH���MO�/WOF;�Z宨¶J1�j"�A��"�Bmy;;���0��0��}�<��WX��Yl�3@\h��`,9�H�WF�)Urx�$����5B%���O�����4��_���e3,��V�.o)�B �nʃ��#�a,n�cqgF&tS�D�H���MO�/WOF;�Z宨¶J1�jn�ţ�Gi��(�V�ܼ������A �׏�����MFi��|��wØ�ߵ���#�!�q`�q��+�e�ZD� �9D^��kGQ��l�4��H��x�d��cɁ#g�k���}?�N�*J������w�����K�Ǒi}3�J��[�
�� ڈ�)�`b�\&A(`#� ��u���'���ߌ[��83�$^Ȟ�]��_�'���ߌ[R)Ms	[��5�(b��g��U-�eO���EWI��X�)Х��=�\2�lFb�A���Q������;e5V�]C���[���?S�*���X:�*��ܟ�8{�g�G�m1�H���W�w��fDИ|��,��9x��i��0aW��➇�~���:�d�p�Pm �5�����	��Uioέ����go�+���}���^���\�}M�/>�96���1@w׬�H����[I��;��A��,W�����K�Ǒi}3�J��۪	�}a?�d���&�ʕ�I���(%�9����p���|���؀.ņ�a�t���EF�w*,�AMX��Qm�"�����{����r�&�O��p��	>;�́�^	�+|~�tݧG �Ŵl�;�w����X�:�{������,�ǰ6y����m��޹���YF��(&�ƫѦ��2�����Vc2�����Vc2�����Vc2�����Vc�]ivc�~�����9�7m����2�E:WK:h��7�������2�����Vc2�����Vc2�����Vc2�����Vc�� ���P�^��P0��JO]�"�?���q.�����'�7I|���;��|B+T�
 �������YY>��9*��gB�Ү�1�f�؇��*����
�?<1@�J�r�f׿�������!N�m��n��&�7a	��������W5�\tCՌV�����,����_,�qo�,ܛ�	��������'�3�$ �#^�Vn���v_�"c�PƐt
׫�J��!��l��[�?2^�9,����_7γҬ�,;r�mR-AF=p�f�[�p.������3�Aq�yo�${U��w�X�|0����p���Φ�"�K�b��Ub�ۙD��׊��s����+8M�?��CGb�% ���+d�@Wێ`�Ӻ��L����~�pP�R���+a�G3�u](⋼�1ވ�'��Ǵϴ`�-2c��ҭ��'���ߌ[��83�$^u������~��j.o�c�\.U1+]2��F�fsxx�rDc�5��ja~��j.o�c�\.U1+]�Ȯ��ߊ�����B}�S�*���X:�*��ܟ�Q���@e�c��1���8}�Ͼ'���ߌ[R)Ms	[��)F��'5x$Q#�&ՠJ�14�~�Xo��0����a�Z)�����z��>x��F�\.��0E'jK���:�^���A~��j.o�c�\.U1+]��:�B�c~���;A���p�����|AW�G�E߻�"��|���kJ��K�}i�e]y]�g�ЄQK4r�n�鬃������-X8l_�m��k�ph���X �����R]Y�/�J3�`��Wa-�>�ٌ��gPǢ R�*�߾�'w��n�Ak����h]f��Q�4���܂Y&#�=å�{��Θ�r�B�,{�H��2���Njr�Ú��k�VX��h=as��9)N�D4�ky��~�ch�B�_�+�)���&���/�����|�*3d��'�W���'hW�S/f��e�WDv�b��h�Ӆ��x��h�6Q�7�0ʓY+��g�$��b܉���5t��v �-�F,�C���� �%�H��,ۙ��*Ը�����
�?<��X̖���Q�$�Wjc��,b�md��4Y0]�Ys2���W�����Es�a�p梯�DΦ��tL��,c3ಙ��%!�t��;�6��X̖�7������qk�	(���f�>Iz�n��VK>�h$G����H��T���+«7SŞ�Ӣ��H M��� C�(��EZ ��07�F��b]�iz�?�d���&�\�S���1!޽�n��3�E��� �g^M�va,�X����_��(K�&?�d���&�h.�M[�̢M8���2	6?�.�
oq��m���k�zm ������YY>{��E1�orǟD�ui9�f?Y�O �iʁ����mm�T�q!Ul]����r�|�G�n=��/ݍSc��6���y�=k^ŧM�m��2�`�W�K�F�����;
�V��nyk��Q@���T~�-���-�\��l��)�>�@#zv�`�"�X����GG�8��F��@���_w���<�U�?��CGb�% ���|�Zqg��B:�N��u��eu��<�'$�x�W¡����O�8HL�N%��**m���F���9�@Zd��`�H�&���1DV�H��~ж� ��%lsσw�kz��Qf=��n�# 0r���q�L�昡��:�C�l�1�ԀU�܄��� MY&#�=åи�]+z�@��.��c`�V�s�]Ҋ��$�R�n��|��KB��0�^��C�k�j{�@�u�g�~�ch�������l#QF�ky��.�"=l�o �<����e�|��ooF�!ݒ�N�PP� *����h��|���kJd��#���G=X��i��?Z4Z��N��b�٥'�E�Jg�S�(��ɒY���ƛLa���Mw G,��L|�:.:]I/���jbPhޛp4�.O�+�AMm?��ˏ8[$0���]��#r��`�3�Q��RU떐V�RDFR7��/
����X?�WGc"�Ee�6;�M��nq����Cf<s0���UY�^����L�Y&Nkj�w�U4~�~��y��Kᷪl?
�A��[�E����7������qk�	(��&JX�=8��������)��[6��e���o!f�	�Ĳ�z��y�J�#z���=����=J8��|��d�p>W< |�;�Ojz�@��Y�rJ�IaF�<��yѡa
qs{a��!��=e��7��5>�l8�c�������yѡa
qs{a�򖒒�����Qs&�1@Җ��{��&^1�ā���} z�U6��0��JO]�"�?���q.�����'����ڇ7��;��|B+T�
 �������YY>��9*��gB�Ү�1�f�؇��*����
�?<1@�J�r��Y*i�~��~���;A���p�����|AW�G�E߻�"��|���kJ��K�}i�e]y]�g�ЄQK4r�n�鬃������-X8l_�m��k�ph���X �����R]Y�/�J3�`��Wa-�>�ٌ��gPǢ R�*�߾�'w��n�Ak����h]f��Q�4���܂Y&#�=å�{��Θ�r�B�,{�H��2���Njr�Ú��k�VX��h=as��9)N�D4�ky��~�ch�B�_�+�)���&���/�����|�*3d��'�W���'hW�S/f��e�WDv�b��h�Ӆ��x��h�6Q�7�0ʓY+��g�$��b܉���5t��v �-�F,�C���� �%�H��,ۙ��*Ը�����
�?<��X̖���Q�$�Wjc��,b�md��4Y0]�Ys2���W�����Es�a�p梯�DΦ��tL��,c3ಙ��%!�t��;�6��X̖�7������qk�	(���f�>Iz�n��VK>�h$G����H��T���+«7SŞ�Ӣ��H M��� C�(��EZ 4b�zvѓ�)s[�3��kd��p'k��o��`��[A+��F�ڪ���B�4����0��Gh1hh�r�qgF���~�v������N�1�� ��2�����Vc��Y7�E ݨ''��*�id����g: k��2�����Vc�cRq>h�3U��8�8�	J鞑t�T�/7H~H=U[�"|�9�GKP�2�����Vc2�����Vc�"��^̹���c@�ȭ�Bס�(ZH4~��2�����Vc2�����Vc�m7���e!�`�(i3��E��Tu!�`�(i3NK8�y ��· ���4!�`�(i3S,5W�+�NEx�̶���}�
�"�!�`�(i3!�`�(i3���w0�!�`�(i3��J���i�X]��w^�=���0;�٣�7�Ƹ.��v�n��v���!�`�(i3!�`�(i3��;I6l��!�`�(i3&��潹!�`�(i3qa�EuK��+���R0L А��&�^C������,"b��\�f_�zH�� �yk�&���LSM��;I6l��!�`�(i3�(]:�z!�`�(i3!�`�(i31������I����!���E��+U�K��D,�Fj��C�ri��X��Pꃅ%��W�c���q�B�ݔ�]<�gk��mZ�+E�Tw�· ���4!�`�(i3h,��3h!�`�(i3!�`�(i3�· ���4m6
�DR�П�� j�L*կ`��%�����-���,���x��
R���eU<�������|[���HHi���~����Us��v�ʻ˸I�d�!�H��· ���4!�`�(i3��J���!�`�(i3!�`�(i3���w0�w<�_֒Hv�[�2���eH�f0���������㗢%����֝�r?4��oH�l��ɸ׼iնԨ��o�`e����ots�SϞ�TsP��)Ԙ+��ｗ��u��?��Q�&{��8�aЉ�O��ڗl��}���^���\�}+���Ã8�4��Q>�9g�M�G�n f�Lu�m9��u�{�C���� �-��4.�B� ��~���4M̍����Q6vmI/5(Q�g�+%f���at�)��d��X��WG ��0/zﴚ�h�X�/����{q�J�)�>�$�>�\�W�ECpa=ja=X����v�� f�Lu�m�
rQa���d��{S�+�AMm?��ˏ8[$0�\�<���+�R'cf���n"��
l�	ACDCx��-��߂��g�K�
��� )H]���؈a����cI��S}H�
rQa��Y]�����V�RDFR7��
rQa��Vf!�q̿	�ZXĒ*C���� �w��wv�G_�:��~����h;�ab���c-(��h�X�/�D"����#CK���L����E`���rw�&�z<a��N� φ��<�6��!�Tc_j��r�.XeN	7J����e�c��n�cqgFz_��q�s|�3�d(]�/{��l��8�[��آ��R��C���� ��#��+��f�iC���(b����Vz�v@��'DRŔ�rUq��ɤa��)gΔc�"F�}�y��Ps_*�GqW�w��fD[�1}[�7HB <��g�^)�+CԼ�xXyN�]<���)Ԙ+��ｗ��u��?��Q�&{��8�a�8�m��;q��Q���F�B�
/Sq��'�E�JgJ�k�ٰ�)�>�$�>�\�W�ECpa=ja=X6UQ�㔩J�k�ٰ��^A��x����
�?<�ޜtW��6j�"Hs�n�g��mW[�Ƶ\���~��c��Rr������Αo��p2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc)_nي3�/?�s�m/C�Ѽ?��Q2�=W�֯�^��N�&��^˻f��)	e�6k$ުm����Y�{'%sAԢ�a\蟔�֔����ߖ�g��o�4��?����DNZ�j׫���?_W�\I��ఽ��`g�5��!08�tw:g�/�6=m�	n� ^�d�#2��0�DQ�L���E�#�K����!�������Χء<\:��{�ϥ3'�Ƞec��	�Ė��<��:-�M��Q<G�^��	#&�^��m^~_cv�;,�Y@��Q�Ę�5xM�����?��9)ٓ���j�2���ع��;H/pH�����qg@ۼ��.s��|� ȼ�׉󾶓:��,�,����|#^�Vn�^ֻ����XP���6��tJ9���BC?T�<o�nïi�JHn��z��r9�3� �����Y~��`�JKݗZ:���'n�^0o����y�]�$�R�n�9j�ʛ�q{�f��a��4�6�t�A��u�#փZ���0��q:i@_�8x<�A!lxM56V��� rJHn��z���G7�����z��>x��F�\.��0�q:i@_�8x<�A!�>߲>���g,�5�Tz3�u,���W'���Xwd�n]N���ۆ7N1ƻ9��[�>�q�E#�UJ�#��Iam�D6�U6q�����20�3p,��ud�M�L�IÙ=�Hz�n1:=��T.?T�K볋���B�|��m|�z��e�i�"�����{���_���wg�|��].��'���XwSn����P>7Xl����]�Jg����-c �ЄW:��2�-4�������A{��JVjN�h�Q�;���T2E�5X�vZ��Bv�~������]�!�����#eH$�DZ� ��o30�@Cd�$�j����"�YVķ�;��h��Jh�]H3=-��7�s|d_!�\�<��z��}�צ:�)7Sx:��7�q��0D?e��{n)��G�D(x��|�e�UTBf����FH^4/��?Ev�~������]�!��_�t&����hx��W����c��a�$Z%�	��J��bZ��b�Bv�~������]�!��j54Z�K�;�q&�<ν_3#ڸZ鎬�������(���}/A;T�c�h���o�8���/���P�ţ���j�b?u |�V���r�^�y4fCx=�a}hU��xz88y�[��8k>6s����]�!�������͋��E��w���8<:XQiҗ�.�����k�fȜ��@��ӟ�x++5xM�����?��9)J Ւ�&�$q��EI]��v�j=U�h�]�vv���E�fZ@IE�U����S8��m�o�&i~G��;ؔa��-)�]��V+m�?��+z�J�k��]��nsמC��_�2��+h���l`�M����޻�F��&���#�{�0;�}���K���sמC��_�2��+h���l`�M���xN�k�ޙߤI�p\�WB��"?�N|I��`�orǟD�uiL${?�����>��yܛ�	��|��	(���zL͊�q���19TH���'�3�$ �#^�Vn�^ֻ����XP��Ȼ4�t=�j�.�/'�����W;5B5Y+� �i7�sp>��8"�@[�f;q�sɈf�=K�:���A0�	}�A�X5��_�G��Gq{�f��a��pP�o�0�CXL�\՚�P�S�bN֕L�����zL͊�q���19TH��wJ�G�����t �JHn��z���G7���_��د��� rJHn��z��^G��OE&� LK�a�]G��wi�bZ��b�Bv�~������]�!��%��rSe�u�heJ��Dv�~������]�!��	Ǹ�y85��r>?�W����/7R�%�T�\ ��
]�T��i}3�J���č�Y���S�)37J*uc�A�L'� |��JM����P�����s�][S���C�ROe�Ё�������Tǥ��| hZ଻|���9�dMbZ鎬�����W-O4�؏�F����U�D�>i�ל3tj�5+����~���U�z	��ߓ]�>k+;��5�k��y׽)N�[SV��˵��W�[4�	�}���^e@��V�i�I��Mֱ�H���� 5+� ��G�|��8��\n$̱̉���ߊ�,�'��.	&'Q����^�[��$*�¹�>D�� ��;����=IEw� e8�~�����0�H��OR�JO��V�RDFR7�h�Qf�����m���t���S�����ۄ؈��k�;4 e8�~���zR���bp;EK�6(��Mށtd؈��k�;4 e8�~���zR���b�W� D���>X[V��kC��8��h�Qf�����m��u&^3X���W��'LC��8��h�Qf�zm_uz�o~��������S&ϊ����֬��g��i�U�T�٥��TZ���dJh2�T�!���j�bKZ(��δ��� ��&�9&�]֞��� �Z���dJh2��9x_�+�O���J�w�@�Va��1_���k�:;5B5Y+��כJϾ�i���@	Q�j���#���«hj)��)s�禖g�đ\e�O���J�w�h��l7^*�Թ��:�l|Ѝ�e%p��\�vş��i�~G��;ؔ/Sy�,v�@�Va��1_���k�:1�*_��h�V�8�]�S�*���X�#Gw6�&(@Y瀉cbp��'@
9��yū�Rm�Ƈ��ݱk4# ����5%JM�T�\ ��k��g��~��j.o�������u3���4XR;�=7�B[&^�D��;�L���9`"����(�6���l ^�V]��}vT�V��|�������c�A�L'M�Kc�Iؙ@�Va��1_���k�:^�V]��}R�wX��pzl��a�V�RDFR7��3w"��R	\{���ͭZ鎬�������(��＂��@ê�Ь%48	>Wٹ!5�j�B�Wǖg3ȓ8���/�P�u���5����������+�ڔGdb�����6�m���d?֙�꧀�s������`�D���>&� �V$��K�Q����
�?<�o[�n�g��R"{�.C�$4�	  Է�/�>EZX��s�oaWZ����m#M�4�B�_�+�)k��G�s3��d�٣��c�A�L'M�Kc�I؆h��l7^*�Թ��:�~�G4PN��g��U-�e%i�8��So����|� ��EX�r���eC��yoZ�P/���dqy�nrm؊(��~����p����
�?<2�,)�<E�����*Tp��:�z���Hhqu!���5�Nn���4L"�#W��xW�Kg!�h���[m���~������a����N���#t����n�~����p�@����9)����K�d���tn�u�$d�I�v`J��U����+=����7�>D�c�lQ@��~�
�KT\�mɍw�B�I:׷�F�20)�_SsJjvCn������Y�
���h$�7�R?�6��%]����	����ѕ��J��<�..�4��?�뭨�fv8���p�lő�4�`�+��t�Y�Ij���0E��@� ��Le��	I���]�HЦ����AS��M4m~�����c-�z��~��D:ǯ3�4���X�E��	�'�J���U�2Gޣסe� <���^[ �1y�,	��"k@:G�	���=�ܾ�y�c��"x�O|?.����!��!����W�������9�xV��	7����G��O�L̍5��+'}����4L"�x��R�>(��F��eTQ�ȋ�V���w	����h _;��i�1�Q�^�� g�!�{5ܛ�	��A����¥��bMݪ��V�����׷eh��S�=�"�56RmHX���!���H���vO�[Jf퀔�������sr���0G3�f�؇��*���Y$���y�z�ۼ��uWU4y5=>F/ġ"���Չ-d��r�b+ӄ�bİ��i+��*�I�GIN�|L9���f�j�M�n����x5=��{t_�sVh�a�|�&�#�E�d���������|��=;��|B����?�IX[��O2 7�,�)�C�BS��g\��ı�ZnZ���qq�c�@,��ڬ�A ������ĎɌ�[9�-�Ҧ�{b�J��@��$L��%��Z��b,�0g���>a��v�<�RohWt�_a�fC��0��:Y����i%��ό�;�LȫԷ�/��Ϥk�;��|B}ø��y�w8#�RC�G�G~��6 ���F��G�z�e�3�ԳN���#t����n���n�".�LV�4�ұ��ݣW�](������(���4,e�b�����E(��6��cd�qS�?�����X)��X�˂��.�����ՒuL"�^�Q�؝yl!��'��K��8�0iT��g*ޘ^��c�R ��`�ϋ��G�m�P�;�V�6�Y�����
�?<���d����V�w˨	R���N-1gΫU *QKE�껐�LqE�����������W�!�LHi�S�������GT�}��K�)��I�-�A`�Mξ�y�j\ؕgD�%u?-/=z��;ٱHp�Rew��i��p&Zc��gc�jv�Тk���aA�h�Ӆ��x�;�琾BT���h�}q���'U�	�YI܁���˺�Q���|�A��^WslxSwP6h���X �.���6y���/\�3�=�7�V��g�$��$����_\�M�9sW�l�l���XU(�a����ؽf���~�ch�B�_�+�)��#��R6�.�iGJ������q�����I)2����x�:��;� ��$L�H�:�z*��y���b?�o�ԛ٩ո����t�:��s8b�.��;��|B���D4�����m#M�4�B�_�+�)?�gγU���q�b�-G���L�{xiR��ٞ��/>x��F�\��Ɲ&�ko��_{[�>x��F�\��R�>�v
�ߴm���bG�~��j.o�c�\.U1+]\Z>�?��"�:�� [ws!<vsH3�3P|�+��?�d���&���gE��Ҝ��z� �;�t%k�Ϧ8k����y���b?�o�ԛ٩ո����t�:��Zcqe�+�;��|B���D4�����m#M�4�B�_�+�)?�gγU���q�b�-G���h�2��>y����,�ǰ�6�Pr�|�1�eP�#�F��v/Br���~�Uioέ����go�+�
���,>�Uioέ����go�+��b�ZhC�#�I�U���2�
PT�4�����uS�b��?,�*+5܊��|�%����0�3p,�;�MRq_�(4���N�3�+�	��o������9Xur�;�LlHő��LA�dWH��Z��Q����Eߧ�� N
�;�p.����������X?f��˚����Z��0/zﴚ�����j���P!3)T�����Y䉪�m#M�4�B�_�+�)���H����m���L[�'%��gXR;�=7�BV��kS똌,0=]^	�&���}D�I4>��z*P�2V�q�Y�*�B�:N=m��
�$�����,�ǰ�6�{���o��5�kd�h1/��	>��< 3LV�4�ұ_ o���5�s�epe�����5�� ��tȈ������<���u��銏�H	��j��|�(�@3l�֮3���O.1��ܐ\5�OYp�V�RDFR7��HwF�E0���'nZ�7�w���"E&��� ��A��ˮ��V�RDFR7��.f.:6�G��O�C�_*�����=֥7$�9D��ty�և�j4̗��W;��"r뾃	��s�G�v}�v*��v�M�����]V�aK�asRF�T��]�w9"x�g�Hz����V_��I"� ������Ewj�,� t!2�B�N���D<����e�cN�Z���dJh2��)���u�̈~����UӇ��ۺ�ۤ�&�L4⭦[fሰ{���Z��0/zﴚ�S��W�Da�P;m̳�}�_�������������W���>��yܛ�	�������,����|#^�Vn��JM���w���BC?T�<o�nïi�� T[��m��U}�	�(��Q|3�@���U@���:��F���Ed8���d&(C�#�7#^�Vn�,��`/[�f;q�s�~�Ԣ��D{5���0�CXL�\՚�P�S�bN��P])Ưbښ��>ܮY"f��g��6.>���m�d�z��*�B�:N=Pp�}��
K����E�<�]�#����$��
��U�_��د��� r�����
L��T�����(f����j�ơ9��&@�E���+$nCe!0�K�r����h�ᮛ�ڥ��!���α�%�����h�f����_�y�&P�i}3�J��h���X ����
�?<=�+�	�;>6���Bi��?Z4Z�SI�(���蜍6���h���R�޳O�
B��$��~a$�BU�౸�������>����,�ǰP���Mt&���tz-��Ű�ȺQ�I~m��Dk��m6[��!N�'�y�G