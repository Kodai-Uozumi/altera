library verilog;
use verilog.vl_types.all;
entity \HCSTRATIX_PRIM_DFFE\ is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end \HCSTRATIX_PRIM_DFFE\;
