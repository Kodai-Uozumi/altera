��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���a?K���J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-���տ��ê�Y�o�:g �C��A�F�7���3�GXS����E@��~���($�J.���
�=W�֯��i@F�5�=h�GD��aC�h�>���SW͟��W��x[����Ȅ�\#+��S��3��3%��׍����}0�st&���\�vūx`��:�֡�\�<7�X�e���V!���IÙ=�H�l��3d�`.�/'�����W;5B5Y+� �i7�sp>�2jL�K�B���.D7�GV��F�-���o��C!T*�q���U����Е� �7Ê7�E�4'���Xw<b��&ɛx�����4�b�k��g���7fj�~���3PS���X��u��(�
t�������2�=�����R�S��q�P ڨ��S���Q�V�ɶ�w�Q�41�&��~�I+����R#e��ds�H��b�^5J_�>�q���U��ȓ�iӚ/��Ϥk�;��|B}ø��y�w���H1��@�	��hN�q;�ǔ10\p c
N1�V&�����O�qTkή�Ádo�dvAg~�rk܀�#��˩���.|��f�ͣŗ�:���+"�9���B�I:׷�F�;�sB*�1v�!���y �谝��X�e�F����To?��m\Ӓ�qܛ�	��]���������ї4�z��pU6�M�S��2�{��΂DЫ�5�E-%Jn��ɧ���7�)a���%}D�����!��g�-��\��OA�=�~�]��d�Y��o�6�֟�Zl��a>���(�WI�;�_�	�t쩖NUD60L����L�Y&#t����n�~����p��l�n�Zl��Ͳ�8�3���!��@HW7��ո\����8�L���9���D�K�X�Re�d���L$�ѸT���C6���$73���'���)w�i����0\p c
N1�V&�����O�qTkή�Ádo�dvAg~�r{m��<�te˩���.|��f�ͣŗ�:���+"�9���B�I:׷�F!���H�v�!���y �谝��X�e�F����To?��m\Ӓ�qܛ�	����%��1����ї4�z��pU6�M�S��2�{��΂DЫ�5�E-%Jn�p�+~� �yKYQs��[�|�F��ˮ�pd�Zз���\��6�R�X�?�I��H���Kn�ǈ�s	\�@0k W�:��S��y9Ez��}��H֞��� �0\��.�g6���@�H	)pH!���5�Nn��XLVt����G��5�On"WW�p��G��8���Y�઩0g���>{@�w�|���*��>
�-�E��{���dʡ��'��gk=���G��yʼɊu�V&��F]�&��yJ�y'��BSz��w����s�%Ƥ�/���d}��[�ƭM��g������Hhqu!���5�Nn���4L"�+�va��2kYD��ʗ��'aOދK-\��$-��Ǡ٥cX@n��U��Y]����o��_�RP�c���
O�KX��ik9�$ C��/}>5��0�x��y�o��ƍgR��r��wėZ�#o�]�ʄ�B��LJ�.N�Ii�,a%��w�J�@R���=�<�^B�R���>_	��$����Mv!���x�5ߧE4��it��ı]`���vuۂ�>����� ��M�W8߸��S�Ȍ�^�l���+:��0	��