// $Id: //dvt/mti/rel/6.4a/src/misc/avm_src/tlm/tlm.svh#1 $
//----------------------------------------------------------------------
//   Copyright 2005-2008 Mentor Graphics Corporation
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----------------------------------------------------------------------

`include "tlm/tlm_ifs.svh"
`include "tlm/tlm_imps.svh"
`include "tlm/avm_ports.svh"
`include "tlm/avm_exports.svh"
`include "tlm/avm_imps.svh"

`include "tlm/tlm_fifos.svh"
`include "tlm/tlm_req_rsp.svh"
