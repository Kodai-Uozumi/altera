// $Id: //dvt/mti/rel/6.4a/src/misc/avm_src/avm_pkg.sv#1 $
//----------------------------------------------------------------------
//   Copyright 2005-2008 Mentor Graphics Corporation
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----------------------------------------------------------------------

package avm_pkg;

//`define AVM_HIERARCHY_DEBUG

`include "utils/avm_version.svh"
`include "reporting/avm_report.svh"
`include "vbase/avm_vbase.svh"
`include "tlm/tlm.svh"
`include "utils/avm_utils.svh"
`include "deprecated/deprecated.svh"

endpackage

