library verilog;
use verilog.vl_types.all;
entity \PRIM_DFFE\ is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end \PRIM_DFFE\;
