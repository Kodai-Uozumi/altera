��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���a?K���J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!��Q�"u�b�c�#3�-{_sh�o�vAg~�r)�t~IV�z�������U��d�ф~����p�1!�΋;Dvn��I�?��]����W���' 㴟��Gn��:6�r���p��VL��*(o���6v3��'Ytp��:;�[���!P��~�|M*Ęj2�B�[�b�x�L(����A.����4��i�%�!�>����O�	
ߗk�J��I�z�]�c���x8��H��Z��{_��iЊW���5ºvB�s~,ptQ���}�L<v��e4�����3dJp��L�8H�@7��G���ږ�3xZVP�Xr�][�@���rah����f�����6�Lq�2,ߏt�Ĵϼ	���6�э�|�����B�3|}s珇�EH%ō���!�X��KȘG%�=p��SjT���O�vq�M�4�H��H�Ǉ&���M�6��v����
#U���:�Q�kv> ���mz�� |��/�Xh��:e[�#�մ�.B;O.��Oz���t ��c���x�6���v���?�֋d���=L���4_�?GQ�.��V��?oj�s�g�7���ϾU};ɀ`;�4���(~�MǓߥp$���"��dZ0o�v�T��^�v!��$0j?�s�����XI�a�f2�[���ٹ���م�uLꏯ<>x�2`�J�É�����d�x����e������k	����UvЅ��Q��j�`�ϋ��GmJ��ɼی(y�3�`�����x���B,'u���/8'�QL&�v��H��2���2�()Ȕ�7� �M��O ��� 1�+�44΄,�H'u$�5�=�7ȸ���<h�<�V�QK�}�Y>�K-85I��ޥ�9���b�j��}�d�܂��Y�kí��K��Gn�*TȷG١��3	[G;�\5�I���(����<��Q��V�ea���}ڌ�� ��1���d�O��{��nrm؊(�p�Y���U�m����]�cS�GN�f�U*�qMC�%`zh��g(>����;�Ӏ�sqS�I)ŢeD��8�>z��4%��짐��R%%F�%��짐�(�N���P�7H����>��E������y�.q�Q�Ҷ�dǙ��
��A|������7�ݒ}dZ0o�vʱ3������6��n��`���n=2�����(å
�A뫰v]uR���C(QGŎ·�K`������l<�Qudw��|@�M���5^s桃��k�Ĳh;�E{-�>�����B�ժ����J�A��\�${i���~�;�m^$��
�/��,�R_cb�
#2y��g??���CM��5�Sz��6�Lq����P/�[�CM��5�Sz֞��� ��� @����eGfFXջ�hʢ!�5�	�����ތsȸ�"rR��(�ٱ�W�I�z�]��&���V�g�TI���P��mgA��k\�����"�9i&�Q0�u���%��짐�(��v�r�]s�ES�T�<L�*-��pޒ�.��P]:�K!��]#5؝��Ү���<Mz�0�4��3�>=���#,J�l�/f#�}N9�h�{JB"���y�#=�h��M���5^s�=�kN�j�����ʂ�)Af@�k�&�厏�c���Z/2�sȸ�"rR�P�΃�F��t�Ძʃ���#_��⋬n��2%0���K+�,x�W��.��贅����c�Ѽ?���FCx��!�`�(i3}C��uo	�l+%��xC��=��:67�,���%�����	����o����ry�TG,���%����(��X> r[B1Y������Fz�<4f/J8�<}�L�Wa��Ĩ4�/T��ê�Kq���a�S�P��3,.x�Ȫ�>�B�HCڰ������c�H���ׇӭ��5�����}Y�e�E*'/	�7.����f��%
�������FP��cC�Ic9S��D�j���r��܊F`��j�.S2ׇӭ��I����d��r�b+ǯ3�4���G2���*�)���K����c�!z�i	'3�=٪	�Z�I�C�8%~��im��ғ�;ab95c�����m��!���"h��1���!im�Ia�|�����>ր 6���%k�����T�:�g??���9��xqw$FD��N�3��뙾�SYO�i�%��!�r����2��O�&cj=�׶�@�$Y�*#�IQ܋�9�2"�!�`�(i3C�A<�Z�̳P�ߙ[qwQ{>�붋"�M~O���ƻo2j�`$|�ku\ad����6�z�
^9�*�l9yt��g4sȸ�"rR��0�&�ͭ���<My�zk98�5��W(��ɗ�s�
>{J�^C���m��o30�@C7��G���ږ�3xZV���)n?����뺨����>=���#Y�J����x���Uͱ�YxM��}�!�`�(i3�Y��nkMM��m�7�TG�>{=�b]!	r��m�z��b6������P��y�#=�h��M���5^s�"��FlXz~�Gy�'W��	]�	���D��ܒ�����[m	���Ʉ �����#(L�̷v2�j!�`�(i3Y�Q3�tY�Dy�-����F>����٭M�3�9��)pZ���b�a�WX3�T?ې!p���.��Щv<�<��hK.���Fz�bˑn�9�Ƅ^�=�]�_Jz���j
a�I���;% ���WyffwA�!�`�(i3�"��kyB��ljrk���Q�4IS88��9/���`���6j��p����]n���Q�lH�K&�\�4�ʈKk�IkY�G�ׇӭ�ц�'T���+Y�������l5,/���=`�*嘌\k%��Ns�$���^O��<!�`�(i3:�8���V����
�?<��2������p����]n��؜v�4�oe��t-߱�~�jf&�~�7��o���̄1��7���Fz��V�52SG���Vd�'�K��{�!�9��&A�����˛q!�`�(i3�LQ&��w+K>�_��c����}��[�P5����N?4Y�1V*���p���h�n�ഛ�r��!�`�(i3:�8���V��yoZ�P/��B���- ��[T� c����}���R�-�촎LQ愥~�����8�/��y:����Fz��ݓ�W���Wtܓ��o5xM�����?��9)7�S�����f���;�[!�`�(i3�LQ&��w,V׋jŀ����Dg�D�M>b�B���Zb���6�z�
^Hj����85I��ޥm�>�
 !�`�(i3:�8���V��A�,�4���/,��YHiJU�4�B��ٴ���j>��	��x<�b�Kf�������1EZYq�A�G�+H�pVl�x�7~�8!��� �)cΝ���g??���CM��5�Sz��*^QP�o4�m�ρ�4��	���z�K�fC���4M=���^���Fz�2Y��kک�@ɤ��ӄ+����<�r<��ou���&�����Q�W0jD��D1��n	�I]��Q*7��0�c�k2�}�sȸ�"rRY�5c�P))�jf&�~�7���p�J�����qZ��B[��_Um-V|S��=�=����ly/Z�Ns�`�ϋ��Gr
6����8X�˞�DG!�`�(i3�N�����>��#����2��cF�a\Y������t潅�����c��R����<Fl�Ř#7⸠z�V[���KdyQ��G�T3$!�`�(i3\zgn�K���&�mN-�07����F��k.J���g�|R��qB$e���)\EH�a���\�����
�Z���R�t�r�B���J{��!�`�(i3q�\E��0\��M��ړ'�al��p�~����p|K�mb�Xm[ �tf�A�����KNJ����� O3�7DY��S#"���vL�
; ��Ң��V�x�3���5»9�����$���y�VJ!���(�a���\�"ߗt��E �_�����	���+��7G�����Ƒ��]��3����%�a� ���k��&3�-��_�s*)F����'n�^0o _xB�I��'���e�D�H%�,��ѝq{�f��aƬ$�n������%�a�z�o���Ή&��?��
�^ֻ����XP�����e�D�� 9
�S^i��zz�=�v{Q���7a["�+�\ e8�~��%�n��UM>�䖜�E]����u���B��C����ЫlJ�k3�7DY��S#"���vL�
; ����-���,���"��y�LN��K��g����R�<�W�C%c�����<�W�C%_Q�ׂړ�;ԍ�D���.��4j�%���.�\�:���M��_(����@N��B�)Y��|K�{ߝ9U�$
���Ԯ�r��z m�������#O!��&M����ቸC�g�vUC+
]/R����3P�d�8!��vp�P}��O��Վ��K�����P��$�͌��=��Bl� �r1� �V}$|~ïSup�xg��j_ R�����"��yd\�q[��LFs�k{�L��9U^�;1��\�v�w�?�b�>޼�\�v�8U#��L����n�P�>�<dspK
�����o�"S+V���n�P�G.�V��f����h����開	����5J�^#9�<��\�v�w�?�b�>޼�\�vř9���=��8���c��wr�4�V�b9���:&�>��s��nt��Qw�c*���l���a��XP���/e��I�c��Lun�1-0b����!p���7x2�v���ãf�$��	�(,�ޚ�Q(��L#�[���#�ZA1��Ο2�K��lJa���B&�m��+Xc\��f{>�,��׌_�ڲ�H�� �h0�Y���P9�B��[p]��J��靤�}O}x[��2��'�.�|IH/Q����R���%�h�x#�L_�ZTI�_	pv�r���SD?��T*�Y�k:D6&_���"��yN��6�J���� 9����Ifp`��<�W�C%c�����<�W�C%����_Wr��;���EWr���G����IÙ=�H
,�L�F��KX��ike.�[(I�n
V~$�<�Q��#Â��&?�y�䃶&f��dx���=E�5ߧE4��k.�C��(�%�d3�����o��j~GM��ANET����|K�{ߝ9U�$
���Ԯ�r��z��@�.��������N�|7M6�e��粉�rԯ��Oi����:���M��A���va�{����2��� ��b�FP&T�p�lq�zL͊�q��C���岎� �1x�it�<��cv̼cf�gr��_.�yE%�m5KWC��D�M٭~��,�����B�R���>_�Z>H@���q�^�ˀX@f�,�"�4�04�jf�9��o�����Pm��k�-<9>��-c������[V���|K�{ߝ��-9����X-�3g#C��/� {��M��_(����@҄���G�۰��{�w��.��W�}��b9���:&�>��s=k�Rm���C����7�uT/]�ߠr��_.�yE���:+�B�R���>_�Z>H@����א��4�04�jf�9��o�����Pm���9o,��~X� ���bWi�l�U�N���%d�-c������5g1hw����:���M��A���va�{����2��� ��b�FP&T�p�lq�zL͊�q��C���岎� �1x�itD���o&MX��WG �����n�O�V�ӯ3k���T۳�͕�𺉓n�O�V
^�<vǚ�#{W��:�?"����a�m����S�1h��$P�	���!���	��n�P�>�<dspK>-[1�p��}K��f<�,=K�F~�?|�[_X��ˆk�=�r���x��Z˻r���5傟����@�C�Vm��+��r�1�L�Xڈ*-�kЄ�0v�a�V��!�Xt<Jd��q�G���oR��5l��5��_8\/HiO���L�~׽Ma(FjxJd���IGD@�F��q:�cU�>�ebÆ����2�݋Sw�����3s�p�����\�v�]�����0F�"8����f���e�$�!�w��2����+FC�ϗ�H6���R3���ԏb$���Ϥk�;��|B}ø��y�w8#�RC�G��mf����*�Jq�mɹd�'��"�y���Oq{�f��aƥ��E\����p�U��o.n���������W�^ֻ����XP���-O/ [р$i��Rp�������О.<�Ȭzn�w�'n�^0o����y�]�\�۟�-?�d���&����{ԕ�h7�{`���������������q�z�e�3�ԳN���#t����n{g�P�mP�+���}b��0UcW�3#��9�e��&Z��i��w��#3������h[�f;q�s;5B5Y+�T�����N���,=3���Z�����Oy�����k2(
�D�lnA:�T��|�BEe��h����KP�i�IÙ=�Hw?pª\��T>>M��A���yoZ�P//c�z�5TֺK�)�͸n.�֫�\_(mѦа8��Q�/�V���3��^_�V-��&'�ɀxm�R��K)�V ���Yq{�f��a�с�'sIP�F@��u�����&��"�t�{�;5B5Y+��mV��5f�͋ v"x�'��9e���RBԄ^�����5�'k���R��K)�|1��Ԕ^ֻ����XP���]��Ϧ_�|�|]�u`e���RBԄ^�����5�'k��y�u�?ƚ�z7���e�����hG�'n�^0o�+#�K>��{�TNJ?�s������X�bvN�c�����g�<s*��"fi	��~��n��C��m֐������e� �m�_�Ҩ�V���
y����R���*����$<���GzL͊�q���sT;��i��м8jqY�F}Yi�n/�rŗ��/�NE��l�q{�f��a�:&�>��s��������=�r{A�9g�M�G�n%{���3���4�+/r��!e����>x�]�V��7��_��T��4N�c� LҪ��9Z��.хxNN�(Ņ�E���V�b�����7!�;ۂ��IÙ=�H3�2�y��+_.��jo�&�˃8���8h6r����@Y�>��E-�=)<k`�m0/���3�[U�Ϋ1�4�A��XP���nl{�T�i�
�u:	�b=�E�7���u�7E�YHOIEW8�՚����+�cc˅RO���t��x���:�#gi�n�i*3��hgN��_����b��nw;�0������XP���R��Q�a`c� LҪ�?"#���18z�QkK�[����U��S����[u@�59��/�O���2t��ӳ�Y�
����.C�M��LG�IÙ=�H�	n�늰�Ȣ�9��>��G0�c���ӳ�Y�
���j�
t<h�76AyW���j�bB����^_�V-��&'�ɀxml�4��H���FÖ<^�q{�f��a�1��]2<�	=T�"E&��� ���yoZ�P/�]=a}��:��e��q�탯;\߰��V���
4�B��ٴ��
Y���}�Zs��as��5�"�r�x×v�XȪ,@�&>�JHn��z���hU��9�OZ+L�ʜ%�j@c�X[�\��!?�d���&�m6
�DR����ʺ�?���5��tR�&@>$!�u�]aL�ɜ���F)��`��z � �o*�vo�-7 �3�V���C��\����V�D���Kb���=���aٚ�o����6��/�6���� 9�������z�Ba����	#���,�+V�RDFR7�Y����0r����
���E�/$z{�Ѿ��h��#���%��#i�~cG���l�4��H���F(�E���/ښ[TJHn��z���YG�s�p$C���<��3�
W��1&&����$j.����.��79=��)^>�b*b  �H�,3�V���C��s�wWIÙ=�H�&8���l�mq���)�:�:O����6#�|ސ�r+�\�(��q@���TL߷�q5�ˉ�Ĭ	4�������x�jk��=y�/�xg�T��-7 �3�V���C�Y�i��x4];ˍH���@E�`�Aovj콙����x�w�.�/P���s ��5Ғ�>S�8�dy��{W(l�4��H���Nx�W�^�U� ���_#8��shƻ9��[�>�q�E#�UJ�#��Iam�D6�U6qW�'n-i�& ܵz��O's;o@�1�9���9M/��:M/������;#���,�+V�RDFR7����_�b狡����
:�
5���4�~wD[����#9Fy7GD@�F��q`E�cvR+G
WW�r>1�C�G��$���
G�|�!<��l�
Q:Õ�)X�J�$�R�n�&�ގ/[ ���=���a�8q�O�4D��Y�Rsۅ�LT�(5�.>ؑ� q�.Pa�wI^+������_�����kf���Jx�]�V�����TI��ԑ�g��@��C$����}��yoZ�P/�i;@��\q.�YF�L�U���;�A+b���5,/�C�
؅��FJ��/��<Ӭ��k�K�ָ������Z�]�O�"�"m;��U��aVN�+�S��t��)k�-ohHeg��|����s�ݺᣄ��C�W#@-�ʳ87��Q7�j�!��>��&pR��a��\�}1�-7 �3�V���C1
&���4];ˍH���@E�`�Aovj콙����x�w�.�/P���s ��5Ғ�>S�8�dy��{W(l�4��H���YM�z}�؅��FJ��/��<Ӭ��k�K�ָ������Z�]�O�"�"m;��U�/��2��'���ߌ[R)Ms	[�����-�2�{�OF8w?pª\��3͗I�+O��P�mO��'��U'j��p�U��o.�14�~�Xo��X���d�٣��c�A�L'b-a��K�aU�uC��v��{�'p#I^R)4�����5�2D�3����hV�:��ڴ�IÙ=�H�&8�����f���V�RDFR7��_���׍)�L�m�M�j`�;�_�2��B�>KJ��|�d��ķQ�xO�����y�� ː��+�w��IQ]~���+�#��V�d����Ԛ�ނ{�!��H�q�&������a
��20��4�|75Ol`V)�l֐�?���q.�����'��Ӥ�nq�IÙ=�H(�Y����>��NJ/��!�#��W+Δ}M��R���q{�f��a�:&�>��s��l�
Q:�A�;#�tױ�1���v�;)����=���aw��@�G��o�������HX�r	�y�L�G�I�[U���z-j>yR�_oݧG �ŴP��CnUc?��d��\�v��wc�}�![=���[](U�C��z��
������y��ٓA�ln�~ �i7�sp>F@��uݧG �ŴP��Cn��Y0C8�}4];ˍH���]&�HF@��uݧG �ŴP��Cnլ���4�L�U���;��n�^-@��M�fIÙ=�H�&8���l�mq���)�:�:O����6#�|ސ�r+�\�(��q�����N�l��u@����-_:�?]#���,�+�B�M�5���&�>,L��]��rň�����r���aM"��N�߄�4�X�)Х��؊�K�H��\�vūx`��:�=���[](U�C��z��0�<��_MÕ�)X�J"��Q����%�8j�<1�9���9MȎ��Mƀ�~'��u��m�.��H�c��1�%�e��G�b�<��]5���\�v��:Y��z��Mm�����X���n�{܎�)�V�H���!n}y���q���U�6�£p�=^�?GQ�.��V��?ojʣ='Xhy����A@�č�Y���S�)37J*uc�A�L'�f?S��ӳ�Y�
�ߪ��wZ�n��[��{_8�Y��=�}�Vݨ�%�fĀ�[�}��|M�9W2�R�E$OK�/�k�IkY�G���VѿZ� f�Lu�ms|d_!�\�<��z��}�0z�cUL���gM�6��A+b��ü~���U��g��U-�ee�@Rv����my$�N��lثl�;c����Ew(�A{d�F��M�9W2�R�E$OK�/�,�	��E"��VѿZ�R���O�C;=B>�ǈ��\�B�ҋX������S8�����)�dB%���O-�#���[�� ��q�%a(􆿳�tP"7��%e��0�UX�Pp42JF�Z��ʝ�>	���n�sӠ�k-q뚸�d���A�Pf�d�:h}�"+�{z �g��\�F�s��M_����
�?<N�Y�N�rb<��z��}�<ͧ�:|C���m9�/����Ew(�9V(;�&���܀�fH�k��v�~������]�!��	Ǹ�y85�V�9cޅU��9؜�%��Wǖg3ȓ8���/�l|�*"k���(ӈ�����w����>��5u�Qkgw��.:� tN���&�%_�DO� �Q�c�,e(}�_3#ڸZ鎬����Ĺ#{���t���@�����%zsӠ�k-q�Wv�A��1=ƌ�F�Y��D�n҃���:'�_���wg�!n}y��p�VU��J}\�=��Ӽ��2��}n	�Z^�t���,2����X�kX������`4�E%v�~������]�!���\B��V��PV�)ڶ�|ceJ�z��eU�e�����T�2���%,J�l�/]��-5L�S|��)����\�6�(�_3#ڸZ鎬����Ĺ#{�������犃�8�Qt�z��eU�e��������Dg��y��tqӴ����s��8�M���e���96��`��Лv�~������]�!���\B��Vjn.����Ϙ�J|�Qz��eU�e��������Dg��y��tqӴ����s��W�u��ó}����w�q��N���OG��_3#ڸZ鎬����Ĺ#{��2A���ϻ$�Zkԑ�]�Jg����-c �ЄW:l�mq���)�:;o�������=VU�����WΓ�Y�mݶ���č�Y���S�)37J*u�,�JL�������d)N�UE�B*�2���u���d���=A�2�S|���f?��� <���eW��H��ě�5/U�rQ��3c/��!`����J��<��z��}�<ͧ�:|C���m9�/s9}B�Ź��ݏ1��𠛕!��L�ވ���ۭNJ?�s�C�,������[GL�����K+I�\�q��N��f�;�>)�~�`�0��|��].��'���Xw�����C��Z_�� ���ѡ�e�LZ\^�e���Eы�`�M7Э���j����H��[n��B��X���WΓ�e'��ǩ����l�u+�v�~������]�!���\B��V�e9O��g��$y�z��eU�e��������Dg��y��tqӴ����s��~�̳o�"�D<�4_�;��	��Z\�i�æu�Q_�}{KS�)37J*u�,�JL�������d͇ :�s��]�Jg����-c �ЄW:l�mq���)�:;o�����p�ǔ|�b�ei�5/U�rQ��3c/��!w=����^<��z��}�<ͧ�:|C���m9�/�!������ݏ1��𠛕!��L�ވ���ۭNJ?�s�C�,����&�2 ���������x��lV��(C6	�YI܁���!n}y��p�VU��J}\�=���T�<�����Z1~�g]�I���B��&���a�%�j@c�}������[
]&M��j���$5�}�����q>�~I� �_3#ڸZ鎬����Ĺ#{���Wl
% ��)ʒ�"��/8'�G~+�3;��\���\ ����@���d}�80�[X�b\g�8>!��J�0N�
���	�Bz���tU`f�g_3#ڸZ鎬�������(���R2�sW��t_-Z��T�\ �͘�f��p�b�z'hۉ)s���Ħ�q��Z1~�g]�I���B�龈4��G	������t4z��w���*#�IQ܋[���,d�܉-`�6�����Up��^��0� �8k>6s����]�!��	Ǹ�y85���~�h�Sü~���U��g��U-�e?�:�Z%�~kE#z��eU�e��������Ӟj��s �׊�8²u�8���=ON��t*�[P{C�#^r�3P���WT�j
�I��w��,�9���������a;�/8'�L
�2�Ot�ky����R� -�*3fN&����6��Ҡ��Nx]<	���rѮ�7]�8k>6s����]�!��	Ǹ�y85�ӓ��������@	Q��"X��[���`m��O���U4��{2l���^���@�d�_C�VJ����̕���(��hG�U�Ƕ�2��c=�_R�0��=��d�����caEyF�8ơ�@IE�U����S8�����)�dl�4��H���t_-Z��T�\ ��Sv[J�1ť�}<�&�/8'�G~+�3;��\���\��k�zph5)�� ��լ���MR�Ӝ�n����։�s/�yf��nͼ<�TD��x��3�]�����_�sL�jGC��w3�Z.��	.�V�~�-�r�e�L�]�തJ��ݏ1��𠛕!��L�ވ���ۭNJ?�s�C�,����Hg8l�6o���m�D��%�r �&M��y��Iۯ�oR��͊�]#���}|��XH�����,>$<�խ5�P���Ыl�W`��b0�^ t�X�	I��'��0�u�}�|8 ձJr�U�;�N���󕏜9���7a	��������W;5B5Y+�Ȩ�� "�6cMH%�]��o+W𩡛�5����`K\P�O����X�e���V!���IÙ=�H�SA���4���BC?T��o+W𩡛�5����`Kˊ�jJ#�}�����О.|��	(���zL͊�q��j\~�vB��.�/'��ɥ���;�N���R���c&;Hb^�G�𿆅6Xsd{>33D!{zL͊�q��e?�y�O��) �YR�TZ@7�s�)��}�OV�
��B���I��'�o�${U��w$Q{mi�q{�f��aơ�x�X��Fj~GM���o��KT-}��"q�ߖQ��,�:Hb^�G�𿆅6Xsd����`\]}��A�"�b���"v�Pkt�����R�u� AT�?�z7����b���p�PWJ��j.Z��$�sӢ�]3�����c��(rKg!�h�0���ͭq#^�VnW�F��F�zL͊�q���	��yW��o�>�9�m��U}�	=�C��a���\�vūx`��:����=�ɤ�c�PƐt
׫�J��;5B5Y+� �i7�sp>��;(�˚�Jz�0���je�Vmf��}S���u�����!F7gZ���'aOދK-\��$-��Ǡ٥L����e]�u�����!�G=X��[���J2~M�G�}�+����+u��)_�������h[�f;q�s;5B5Y+��2tCH����,=3���Z�����Oy�����k2(
�D�lnA:��2Y���g��v�x��� T2��zL͊�q��T��Db
�o݆g���V�RDFR7�z�k�Bm��y?h�g&2�(K��ӿ����
Ym�����俧:zvkZ���6�� ���S%�eL)�1��bMI�����^ֻ����XP������a��l)�1��b�:���rw��)^G�<�zL͊�q��j�[���'�`Uv��*(l��(�~�������k��wh0%���dҺt��J��#Y��Ѽ�\�v���'ٍ&�cx�T �SNÕ�*lSf�IO�Ÿ��t+���/��2��w�\	_S>�xH���B){a�N*��XP������<����Dg��y��tq����A��(o�FP�١�&Y��V�$�Ƣ�/몱z���ۀm{�+{*N,=����/�C�ټ�)_����q{�7��)��}�OV9�a��j=IÙ=�H�Z�f�-�i��м8jqY���SހS�ɋ��ă�s;�B�;5B5Y+� �i7�sp>X�X�'��m�Ȕ�1���c]���;�"�!1�U��`__��g��|���y�~��ۢ��9��i��^z\�{�TDHu@�w_���(8@���c]���;�P�����ʜ耚ҵԼ�\�vŠ�B��닶	��};J9��1@��
�b*���t��祣��G=X��1x<�`�Oķ{y(����5�'n�^0o�+#��D�T̻6��v���[�SӠ� �9g�M�G�nʏ�(Z�ϯD�x�&��?GQ�.�b��, �k��G=X��7Sx:��yi����S(���S~���)_�T��|�BE���`B�,�'`��zL͊�q��G�D�� ��|��vt۱���[U�˵�a��݌9�;����[�4-�By��R�i&�V����Sv� O`S�KW�*�	S��ڪ�����$�R�n�m.�>"�RX+�/�o�IÙ=�Hw?pª\��l�mq���)�:��j8HQ��e�z���V�RDFR7������`��I�t?�_��B�e�D�*�Y�p�Yч���Ҟ�+�����ڪ����y��{W(l�4��H��?d�����x�]�V���(c���^�����ܐ�!V��>�%�yZM�����k+�ZG��=�`#7l�;����C���1&&���O�耟օ�[[_rvNH��i�@^g��݀�����oQd�#�e��Fr	�&�L4⭦�����.����w�'n�^0o.�g��R��$���'��j�F7�D�>��؆&,��xA�x�P�~�o��	d��p����ct��~wD[��1O ��tF��XP������<����Dg��y��tq��*��|`�|R�:
��\|��eA&��9��k!�7�D�>����B�Vί��C���1&&����7��߽�-7 �3�V���C�Y�i��x4];ˍH���@E�`�Aovj콙����x�w�.�/P���s ��5�A\���ޯL�U���;�A+b��]j����؅��FJ��/��<Ӭ��k�K�ָ������Z�]�O�"�"m;��U,��BpLÕ�)X�J�$�R�n)��k��U���=���a�8q�O�4D��Y�Rsۅ�LT�(5�.>ؑ� q�.Pa�wW�'n-i�& ܵz���K�ޛzp1�9���9M/��:M/������;#���,�+V�RDFR7����_�b�W󛂀3��-7 �3�V���C�4t����4];ˍH���@E�`�Aovj콙����x�w�.�/P���s ��5�A\���ޯL�U���;�A+b��@=��˓4 ؅��FJ��/��<Ӭ��k�K�ָ������Z�]�O�"�"m;��U,��BpLÕ�)X�J�$�R�n!�OE"X.9���=���a�8q�O�4D��Y�Rsۅ�LT�(5�.>ؑ� q�.Pa�wW�'n-i�& ܵz�rApV�q5�1�9���9M/��:M/������;#���,�+V�RDFR7����_�b�W󛂀3��-7 �3�V���C1
&���4];ˍH���@E�`�Aovj콙����x�w�.�/P���s ��5�A\���ޯL�U���;�A+b�����1��GD@�F��q`E�cvR+G
WW�r>1�C�G��$���
G�|�!<��ڪ������Rm�Ƈ��ݱk4# {pp�����Z�>)��.�g��3�;Y[�i��g/70��� ��E3�]��a A�����>x��F�\Sx�lޞ��rs�i���l?����b��.TpRWl0E���n���7�Ix���Ӻ��L����~�pJHn��z���hU��9&�P챘>,L�ll���(��i�y���c]���;�`�o���PPV��ķ���4];ˍH�c�X��w/Q5���wO�
e�&rV�A���;'Е�k��Dp��";#�lT&A.�������$zz���Gw�� �*b�A䊙=�`�o���]�,/�PM��s�f�3Y���� �i7�sp>5��aF�~�c,�$��1�2>�1$��_w���<�UJHn��z��r9�3,��BpL�A�;#�tױ�1���v�;)����=���aw��@�G���?��z�|걉�BI�j�?x����6�� ���S%�eL)6��9��xx�rDc�ቩW<$ԣ�������T�����N5��aF�~B%���O-�#���[�vE�s�
;'�h$x(�'n�^0o����y�]=���[](U�C��z����7��j�5�i�6T�t�U� ���_����)|f��V�b�1�RR�,�*Ǚ62�4�ͻs�	Õ�)X�J"��Q����j{n�}�R �i7�sp>5��aF�~B%���O-�#���[�"yd��N�}�g,�5�TzS�@/{�&q{�f��a�:&�>��s��ڪ����ݧG �ŴP��Cn^�\���ĉq�p�F><1���ĈL���U� ���_Y�B~�����ڪ����ݧG �ŴP��Cn��g�K�
��$�~ȣ���XP������/D�!"O�p � ���X���n���Z[�ae!0�K�_3#ڸZ鎬�����r44���Y��sx��KK��~4"<��q��P�Zj����(���e����{l�f|��rs�i��=29��aS��na9��Wǖg3ȓ8���/�l|�*"k���(ӈ�����w���{ET�\�h}�"+�{z�)�� �r*Q�%ꐑ�������
��'\�|^��+��_3#ڸZ鎬�������(���0ե�^ag��v�x���owђN�~��ł�!r�dN�<@Iv��nt=:��?���j�B�ݔ�]<�8��0�uM�CA�j�rb���jO��%17�}�w!�c��Bmy;;���0��0��}���*�.Z鎬�������(���d�O�'@i1�RR�,�*Ǚ62��Wǖg3ȓ8���/�l|�*"k���(ӈ����P�`9M$z����fI�j�?x��u9� ȫ^�F3�\�՞&�3�%� \��,�f��ˏ8[$0��g��4��ҋX����L$�����/�{��U��+[+pg&1�����Z�^�\9�����`��fH�k��v�~������]�!��	Ǹ�y85�V�9cޅU��9؜�%��Wǖg3ȓ8���/�l|�*"k���(ӈ�����w����>��5u�Qkgw��.:� tN���&�%_�DOօP0��p���Z۳
0.v�~������]�!���\B��V��HR�gD걉�BI�j�?x���;�Ӏ�b!��u���^d�?8�_���׍)��7�l�:Q��Ig`i�ҋX����L$�����/�{��U��+u�e�+����nU��\�x�/8'��6�m�-~)Ji?N�l�|��].��'���Xw�����C��ED0 � ���ѡ�e�LZ\^ �@'�ZX-\���j�ɡgJ�ت��4/w��+��+r��B��+��|��].��'���Xw�����C�Df�vz�B��{��쭑/8'�G~+�3;��\���\��k�zph5)�� ���;"Q�R�Ҥ;�\�e��`��Лv�~������]�!���\B��Vjn.����Ϙ�J|�Qz��eU�e��������Dg��y��tqӴ����s��W�u��ó}����w�q��N���3�Mo��v�~������]�!���\B��V��HR�gDhx�b縇�,2�����^���@�d�_C�VJ����̕���(��hG�U�Ƕ�2��c=�_RL�2�r�� �w�-}�<��z��}�<ͧ�:|C���m9�/xuK)��d ���ѡ�e�LZ\^�e���Eы�`�M7Э���j��S,;V��bs��OmG��Y�Ȅ�f�;�>)ʣ����I�|��].��'���Xw�����C�F��Fy�. ���ѡ�e�LZ\^�e���Eы�`�M7Э���j�ҹ���9���ϸ�Q�E�"�D<�|��k<�h"r����Mz��;��ҋX����L$�����/�{��U��+`�p�JJ܇�,2�����^���@�d�_C�VJ����̕���(��hw���B���ei�g�������c�,�[`��;��Ps�\�!n}y��p�VU��J}\�=���܃��S�KZ1~�g]�I���B��&���a�%�j@c�rn7Zմ#&;R���_H�6��q��N�e'��ǩ��b�N~�+_3#ڸZ鎬����Ĺ#{����Aدo�zea���||��/8'�G~+�3;��\���\��k�zph5)�� �T�5B���"�D<�|��k<���I�}j����CX�ҋX����L$�����/�{��U��+�I_�=0<��,2�����^���@�d�_C�VJ����̕���(��h��f�<�K6���x��Bm�5
��	�YI܁���!n}y��p�VU��J}\�=���T�<�����Z1~�g]�I���B��&���a�%�j@c�}������[
]&M��j���$5�}�����qwZ K�Ϋ�v�~������]�!���\B��V�e9O���/�\� Dz��eU�e��������Dg��y��tq�2QcV�fV_�mD�ʮ�)���I�N+?^�Fu��<�=��ͬ8�.��č�Y���S�)37J*uc�A�L'�f?S��|�b�@a(􆿳�tP"7��%e��0�U8����p��.?-��o@�e6qR5L�/8'�L
�2�Ot����F�2�v����o/�;�����=f��9c����3��q|��l_�؆�PĔ�5������:�TD���rs�i��=29��a\e�L����owђN�~��&�t�)G9��f1�p!!v*!��u���d�Ӵ���)�jj���|}��3�G��T���93�����wdU�'���띚<�7�6�vg;Je'���Xw�}�瓀�p!!v*!��u���d�Ӵ���)�jj���|}�,J�l�/m�	%�o@U���ry����{D��9]��6�vg;Je'���Xwd�n]Nٙ�mA��ּ��kV���g��U-�e�G:u����# �LW�z��eU�e��������Dg��y��tqӴ����s���w�u1�	�q��N���'\�|^�^�h5���WT�j
�I��w��,c�A�L'�f?S�$�R�n�Wǖg3ȓ8���/���.-�wW��,��e�LZ\^�e���Eы�`�M7Э���j��a:��8<�I�3��
ip@ Iw"���։�s/�yf��nͼ<�TD��x��3�]�����_�sL�jGC��w3�Z.��	.�V�~�-�r�e�L�]�തJ��ݏ1��𠛕!��L�ވ���ۭNJ?�s�C�,����Hg8l�6o���m�D�P�'�h�&�F����U��~T���ٿ�n�P�������h=��
IǬ�{��&�R1˚�Jz�0���je�Vm@�Ɇ�hq��P$��j���}���_x:�YY������8�
Hgؙ��0���2�C���(��
�����Y��/0'~�����_L�{v�B��=Z�˞���7�$�G�j/����X�e����j�J?J��׍����W��s�/Q�-�=p���BC?T�٥����E�?��nc�;È:�-1���{0Yaf�fL�!ȭ�n�h�е������ɧ���7�)a���%}D�����!��g�-��\��OA�=�~�]��d�Y��o�6�֟�Zl��a>���(�WI�;�_�	�t쩖NUD60L����L�Y&#t����n�~����p��l�n�Zl��Ͳ�8�3���!��@HW7��ո\����8�L���9���D�K�X�Re�d���L$�ѸT���C6���$73���'���)w�i����0\p c
N1�V&�����O�qTkή�Ádo�dvAg~�r{m��<�te˩���.|��f�ͣŗ�:���+"�9���B�I:׷�F!���H�v�!���y �谝��X�e�F����To?��m\Ӓ�qܛ�	����%��1����ї4�z��pU6�M�S��2�{��΂Pkt����:a���%�8���p�lő�4�`�+��t�Y�Ij���0E��@� ��Le��	I���]�HЦ��ښ"�C::����������c-�z��~��D:<^��`Y�F�����I��<�|��F+��4���LT K���Db�J��@��$L��%��Z��b,�A�zP��`�� ��D�F]�&��yJ��o�y��e����#"!��4DE'|�&�#�E�d��������y��Ld_&�Q���˛:���,�.ǯ3�4������$�A%q�
�$-���$73���'���))~�� ��-[�v:v�o���+����7X��U�?	r��Z��|�;oYu��>��
��������0��8Xz	fo&�Kh��+�'Pkt���ڙ:t�$Ҥ<��oR���7�m��=�EV�\>������������g�R�"������h[�f;q�s\���L>�Mê�[���#��r�qi�á[�{Ut��\���L>�l�4��H����y�j\k��
3����&��B�cm�Ϯ�Y�����Q����G���#��r�)�1��b�:���rww�u���hil�C���S�V���JH�q��hil�C��v��NrY��8:q.Y��Y�����dҺt�ֹ@���ew������|Dm���v�@a��R\���L>�y�u�?ƚ�z7���e�*m��i�����q{�7��)��}�OVZD�LCZ������ޙ�h��b��1��ڪ����o�${U��w������y���=Iza�y�ܳ��8��4�+/r��!e����>�R�1���4�+/r�pd N^g�2Y���p.������$���{��x��<�����`B�3�!=�ʆqi�á[�l��%������<!�=X�f`�g�W���?�y)����q�/L�U���;�A+b��$���qP�́	P6���y��{W(l�4��H��y�=k^ŧM��ڪ�����$�R�n,�	�X��?�Z
AA��!�=X�p.�����4���Z�)Љ9�������C������_�����Tf�s����)^>�b*b  �H�,3�V���C�7
W��;I^+������_����x4cg��bC���>SELÕ�)X�J�$�R�n���;h<d�
5���4�~wD[��3B��r]�q�D�?�e�& ܵz��<;��إf��ڪ����y��{W(l�4��H��װ��:��o�-7 �3�V���C
�Y���y��aVN�+�S��t��)5����F��\���L>�L�U���;�A+b�햅,��hI^+������_�����\��5�D���>SELÕ�)X�J�$�R�n'���
5���4�~wD[����s�u�q�D�?�e�& ܵz��'~ı|���ڪ����y��{W(l�4��H����V��5e��-7 �3�V���C��Vx*Ж�aVN�+�S��t��)k�-ohHe\���L>�L�U���;�A+b��x��H� �I^+������_�������T��q���>SELÕ�)X�J�$�R�n�]Ke��Kr�
5���4�~wD[���`hiz�VF-|��S��t��)�4���y��e$ׄ� A�����>x��F�\.��0.�l����14�~�Xo��0���l�2q;H�-���m�̳~��j.o���y(�dǌ��E����~��j.o�{���Ʋ��\|��Ea+a�G3�u]����ynɘ�(t�	��i|Stߛ��ȉ26���V�b�����7!�?��CGl`V)�l֐��y�j\��V�b���E9k��-��g<�V1G��_q=l`V)�l֐r��F�$���qP����q�/�`�o���]�,/�PM��s�f�,}%@��`�o���]�,/�PM��s�fն@�%/�w�a�E3t��,B���DrjU�qf���L00�ݭ�<l���@F�K�D��j��'���MIM�աRC U�<��d�q����NJ/��!�#��W+Δ}M��R������q�/i�2��t���������U�~�=]j����1���8�D���kw�т�s���?�������r���aM"����*������+�p�U�C��z����(�~e���(��ʎm�.��H�c��1���ܫjc1��y���:Ḿ	P6���ݧG �ŴP��CnT�c�HfB1c��s�f�=���[](U�C��z����7��j�5Iߙ2�r�)6��9��xx�rDcѴ��B�66�ȷ�	�������;e5V�]C��m͡r��b  �H�,!ԱX�|��\/h��J'��+�p�U�C��z���`�t�yU_� 4P/�W��[�&�pR<�K����q�/B%���O-�#���[�"yd��N�}�g,�5�TzS�@/{�&́	P6���ݧG �ŴP��Cn**�8����>x��F�\�D�E�
���ڪ����ݧG �ŴP��Cn^�\���ĉq�p�F><1���b��#J�/�)6��9��xx�rDc�E|s���J���l���8��!����KsFԙ�0s���?�������r���aM"�������4�1�1�d�$�B%���O-�#���[���)gΔc���T�����(f���5�r*Iީ탾�Q�0�	���Z��zOM���&xg���'UȨ������zG�O�] ���|��&V���2}���'\�|^��+��r����h�Y5̹�����*��Z��Y�N�r�mrۤG�#r�\���(.6���.�4R���O�C;=B>���	����օP0��p���Z۳
0.��v·��H���MO�/�V|G/��0/zﴚƾ>�Cbe�|���A�Cm���Â��㯈h���X �:�}}�I�龔�Π�h���X �/i��r��KI�;����!��ZB4���j���\�6�(���P��
��e�Jh�m��˲��8��1_t�!"�R6�.�ap7�L�(�+�UC�3|�&�Z�oO�q����#���o"��\u��tc�,�[`�z��s@CrH��i�׻[%�lM0��Uxslޜ�c�,�[`�9+��d@�rH��i�׻����{�T��Uxslޜ�c�,�[`��;��Ps�\�7�gI�����ǈݻy<�u��c��f�;�>)ʡ2F�������ߗ�H���3c/��!�Iz��޹��f�;�>)��5�g���ߗ�H���3c/��!��)���Q;�m��H���+u��oE��cFl����h4c��+��#�v�ͬ8�.�h���X ���.#P���������!��ZB�m!��,n�8c.K���!��ZB�(����;ry����{D��9]�~ж� ��%�L�t��n��@�7 f�Lu�m�B�>�9���6�����։�s/�W�J�=�<��։�s/��Wjc��,b�md��t�'wh��� �:&�L~΄gO�3f��*�����&:n�Zp��}K��f<�,=K�F~�?|�[_X��ˆk�=�r���x�i��p�7��Z鎬����@�Q�2�s�JFAa�ߖ�g��o�4��?����DNZ�j׫���?_W�\I��ఽ��`g�M��n\��f[��<j��y�~/r�I��
����&�ɬ� VU+I�©�l|�T�.5b�2��g<3NB����Zjj�.�)7Gx���� ����ޙB!72,w���~�?|�[_	E���=�[4�l6�Pr"?uK!�����
; ���N�N��uZoO�=����'�ނ�ebÆ���p��'ﱑ�c���o�t+����ebÆ���°��W*��׉󾶓:�7�:3w��Ϥk�;��|B}ø��y�w8#�RC�G��mf����*�Jq�mɹd�'��"�y���Oq{�f��aƥ��E\����p�U��o.n���������W�^ֻ����XP���-O/ [р$i��Rp�������О.<�Ȭzn�w�'n�^0o����y�]�\�۟�-?�d���&����{ԕ�h7�{`���������������q�z�e�3�ԳN���#t����n{g�P�mP�+���}b��0UcW�3#��9�e��&Z��i��w��#3������h[�f;q�s;5B5Y+��2tCH����,=3���Z�����Oy�����k2(
�D�lnA:�T��|�BEe��h����KP�i�IÙ=�Hѩ�i�T>>M��A���yoZ�P//c�z�5TֺK�)�͑�d�¶�F���zP��O�O��1��j�P,Q'�_��z�Ӷ�;r�x�9؜�%���5��8�t��\�v�)��+�}�k��
3�����i�V�oE^M�<JHn��z��Wђ�c<�ҵco�SߣǬF��q�~����p ���Oj�r��;r�x�9؜�%��n�F�|q{�f��a�����vo��9ʥ�0
%<d��2�d �~����p ���Oj�r�p�U��o.�ERo�A�J�:�#5��]�W�)g��IÙ=�H�&8���l�mq���)�:x�fr������R�f7�o�u�/1<@fA3c�5�!�7D{�+{*N,=����/�C�ټ�)_�����[u@�59���^ֻ����XP����ˀTdH�gX�(��
���~xCs('w~U���"q���!]���pxJHn��z���hU��9��9��K��Z��	�6�&�����h7�mEox�>�tzo��4];ˍH���Vch�V��\��2U\���\��鎣Z!�X`��_/
������n�,e����+8M�^ֻ����XP������&,5�= ����8������iיf���L00�ݭ�<l�W�U3�hy3zL͊�q�� Ky��:~'���#L�Ѱ�J6���z��K{�̎��#4����ٵf�
]�if#�}N9�h���q �hx��W�B*S�n%w]Ů�٦��l_�F��qi�á[�6���l �^ֻ����XP������4�ؤ���~��V�RDFR7���U�0��S2/GYF��/�XD����@��-m��զR�Þ~C[ w��մ�7}T��|�BED0r➜~y��Y�I��q{�f��a��4�6�t�H�2Da���`�M7Э7l��A���;��|B�X�9�[.�5t��v���R=�;@Х |�8�}7E��O��O
+@~`��)�j�����x�d��I^+������_�����������ĈL���U� ���_Y�B~�����sr���oJo�w���#�lT&A.����4mB�2�1��o�ʳ87��Q7�j�!��>��~�h/����'5��WPu/����Ӡ�w��2D�A"m�/��F��PvF��oE��A+b����ʘ��"l�;�w���q{�f��a��4�6�t�|��+�Fy����N��jk��=y�/>!R3Gb�ǮAi�.�C������C������_����b�o�H�zL͊�q�� Ky��:~d�_C�VJ����̕��W���x��%	#���H�	�q�@S%�����1&&��=ql��.�C$����}��yoZ�P/$zoRؗEII^+������_����x4cg��bCx�]�V�����TI��ԑ�g��@��C$����}��yoZ�P/�i;@��\q.�YF�L�U���;�A+b��]j����؅��FJ��/��<Ӭ��k�K�ָ������Z�]�O�"�"m;��U��aVN�+�S��t��)������Bg��|����s�ݺᣄ��C�W#@-�ʳ87��Q7�j�!��>��&pR��a��\�}1�-7 �3�V���CaP�M���4];ˍH���@E�`�Aovj콙����x�w�.�/P���s ��5Ғ�>S�8�dy��{W(l�4��H���3�C�]�U� ���_#8��shƻ9��[�>�q�E#�UJ�#��Iam�D6�U6qW�'n-i�& ܵz��f�^q O1�9���9M/��:M/������;#���,�+V�RDFR7����_�b狡����
:�
5���4�~wD[��!^��<GD@�F��q`E�cvR+G
WW�r>1�C�G��$���
G�|�!<��l�
Q:Õ�)X�J�$�R�n��X�\�����=���a�8q�O�4D��Y�Rsۅ�LT�(5�.>ؑ� q�.Pa�wI^+������_�������T��qx�]�V�����TI��ԑ�g��@��C$����}��yoZ�P/�i;@��\q.�YF�L�U���;�A+b�����1��GD@�F��q`E�cvR+G
WW�r>1�C�G��$���
G�|�!<�p�U��o.�14�~�Xo��0���p�49k`���&��J�G�D�� ��+G�މ?�3LB�A5�z�}��ƍ���<$���Rm�Ƈ�hʨ}s���ﻋ-�����S8�E�qVf>��6z�`ئ���4L"�k��ci6�l5v�I�D���t�:�S��*~�nzL͊�q�� Ky��:~^� P���&����3{K�貟��N�k�n�,e�P���P����ӑ7�\�V�D���Kb���=���a�X$���w/Q5���wO�
eԥtC��R��V�b���E9k�v��=ݏ�2X8A�Q+����\�vūx`��:�ެ\�+f$߈�vJVt�l�褻�sv���-q]IÙ=�H(�Y����>я\IK�U�RR�%�����}�GD@�F��q�b���V̬���	p�ϴrׄ�ʅ)��~�$G�F�ǯ�l_�F��)6��9��xx�rDc�ቩW<$ԣ�������T�����NF@��uݧG �ŴP��CnT�c�HfB�{���<3zL͊�q������)6��9��xx�rDcѴ��B�66���E���rֈR�-a���O��)6��9��xx�rDc�;��k�Q�C�������P'Q^�	�����\�vūx`��:�=���[](U�C��z����Ջ�/Cp�14�~�Xo��0���$��c����zL͊�q������)6��9��xx�rDc�E|s���J���l���8��!���ķ���4];ˍH��Ȏ�r�x����ה�����;e5V�]C����gg˃xgף�d��zL͊�q���|��3%-�"����}��Ѡ�i�L샾�Q�0�	�A�����<��z��}�צ:�)�]7�˺�9/���`���6jx]<	���heJ��D_3#ڸZ鎬�������(���f�,���Kx�]}�a(􆿳�tP"7��%e��0�U8����p��c���6�
��\=����`3���j�w M��b�%���ؼI�־�2�h�ˏ8[$0���V�2K2S�)37J*uc�A�L'�f?S�$�R�n�Wǖg3ȓ8���/�l|�*"k���(ӈ�����w��2+i�27�yӘ�즤��`3���j�w M��b�M%:p^�vi9� 6*�\�RӲ�I�j�?x��&�nw���]�!��	Ǹ�y85��92�EZ;�����r���aM"���t_-Z��T�\ �͘�f��p�b�z'hۉ)�$q&PbO/c<�2�}�K� Y�tH������)�� Ċ}�MGQ�,�'��.	�&�3�%� 9�	н
o/5t��v�č�Y���S�)37J*u�,�JL�������d2+i�27�e����8����E�2���R/%�|��].��'���Xwd�n]N�m� ��>aQ����G��owђN�~��ł�!r�dN�<@Iv��nt=:��?���j���^�"B{j��&z�D� �i���K�3�"��H���MO�/�����!n}y��p�VU��J)��� �WǍ��?
K� Y���m(s�'"��~Ǣ��t�����y5F�x9xx�	^���龔�Π��č�Y���S�)37J*u�,�JL�������d�q�K�Z�� ���ѡ�e�LZ\^�G�ZN,`��B�ip��{l�f|��:2QYeƈ �-u���k�� ��3d�B*�2���u���d��H������TH-��K�,I�@�"|lKZϖ�L���O'����u9j1�f<��z��}�<ͧ�:|C���m9�/��M�B�J��B*�2���u���d���=A�2�S|���f?��� <H�븑���@Av61u�O�ʹ���B�ip��{l�f|��:2QYeƈ �-u���kS̅��|�B*�2���u���d���=A�2�S|���f?��� <�?W�&����t��!`(HYz�>��A��\35������:<��z��}�<ͧ�:|C���m9�/�T�;��Z1~�g]�I���B��&���a�%�j@c�rn7Zմ#&�ٸ;nR��v��ҍ�!I���Kw�g�P_���!n}y��p�VU��J}\�=��ӿ�y��(e��� �2^�z��eU�e��������Dg��y��tqӴ����s��=���*� ��WΓ�e'��ǩ���KT��I_3#ڸZ鎬����Ĺ#{����y"�'�ea���||��/8'�G~+�3;��\���\��k�zph5)�� ������0����N��� 	�� h"r����Mz��;��ҋX����L$�����/�{��U��+`�p�JJ܇�,2�����^���@�d�_C�VJ����̕���(��hw���B���ei�5/U�rQ��3c/��!lG�g�@��{l�f|��:2QYeƈ �-u���k1q7{�q�B*�2���u���d���=A�2�S|���f?��� <�"��=aet�V܉i��d�=i"}�۞h�G��+^zO��!n}y��p�VU��J}\�=�������X��Z1~�g]�I���B��&���a�%�j@c�rn7Zմ#&9�� :ܝ}���D]��WΓ�e'��ǩ��>F�q�u�>_3#ڸZ鎬����Ĺ#{���x���ea���||��/8'�G~+�3;��\���\��k�zph5)�� �K}�V�h�;"�D<�n�����[�č�Y���S�)37J*u�,�JL�������d�`�%�]�]�Jg����-c �ЄW:l�mq���)�:�ۇT�0��e�zt�z��Al�q�.y �vd�7P��T�<��z��}�<ͧ�:|C���m9�/��W�f��ݏ1��𠛕!��L�ވ���ۭNJ?�s����W����U���d�^���|xV��󉀏�UEs�@�V�Ca��x�jT%q�#�<��z��}�0z�cUL���gM�6�5^��7��ߪ��wZ�n��[��{_8�Y��=�}�VݨG}�tL�x�N=�0��]�Jg����-c �ЄW:qBbr�a��\�"ߗt� ��wg|,���%�̈́T�٥��T� �73w���(���5������:�TD���rs�i��=29��a\e�L����owђN�~��&�t�)G9��f1�p!!v*!��u���d�Ӵ���)�jj���|}��3�G��T���93�����}��8���n��9�n��(�
t�ژq���U���(�M�D�bó=��!��L����犷��r��\Uo"S���B���Ԕjݭ#��2�cv�ϮT�� ��u���}��Y!��TD���rs�i��=29��aS��na9��Wǖg3ȓ8���/���.-�wW��,��e�LZ\^�e���Eы�`�M7Э���j��a:��8<�I�3��
ip@
�L2�Y5̹���^��0� ��6�vg;Je'���Xwd�n]Nَ+vW.�e��h����ߪ��w��ѫ���;�T�;�톇D�bó=��!��L�ވ���ۭNJ?�s�C�,����Hg8l�6o���m�D���3'�L�B�����8k>6s����]�!���)��ɖ�S7⸠z�V[�-jɸ����g����R.�C<�I��ZA���e6qR5L�/8'�G~+�3;��\���\��k�zph5)�� ��լ���MR�����æt������́����H�����Ыlۯ6+�Qq�������R(��z�j�;9�e��ȭ�n�h�oʌjtҫ��/a��w%^ t�X�	I��'��0�u�}�|8 ձJr�U��%�a�"�a�T�r�k�y'��a���4�a@�q{�f��aơ�x�X��Fj~GM���o��KT-}������f��d��]���לo�	�&��$�B�I:׷�F׫�J��q{�f��aƨ:bN�t�ɹd�'��"������JI��'��'�3�$ �#^�Vn�^ֻ����XP���8TJ�����[T�)��������JI��'�@���U@���:��F���V!���IÙ=�Hٍ���]c�PƐt
�2c�'z4�<YG��?b��0UcW��*��w
j$�ëVq�~�I��'�������@��Zdf;5B5Y+� �i7�sp>1�*_��h$)��)��F��arb��@�zL͊�q��K��e�m��/=3\H��^#�6����g׺bH�q{�f��a�P9b����%�a�j��CK]��n��>7n�֕L�����zL͊�q�� �^�ߏ'E/=3\H��^#�6����Q��\�ݔ^ֻ����XP���b���D|ۂ��jǱ��*|V��rP��b]���'n�^0oˁ��6u][I��'���������`C��^ֻ����XP��Ȭ�8�4)r�|ۂ��jǱ��^J���F_D:�	��Z����v��6��XP���9���D_Jx��W@h�l��_@u{� ��%�a�`��]�E$�x7,�V ;5B5Y+�K�:��mA���h{�'�h�
�9[�5����`K��D�	a������T�|��{�r�\	��rR�;5B5Y+�^P/��Ij 4<��`lH[�k�y'��a���4�a@�c�w�V��R���c&;S��na9����:�?i�����\�v��Z|L$ŕ� �GQ�V.�g�.�m�.��H�c��1���ܫjc1��y���:Mb��f����5����`K���\�]\���e�Q8-�^\JHn��z��nw=����o�F�\���e�Q��ݝ� �zI��'�LOi�xg�|��Q;��I�^ֻ�����=�F-�Hb^�G�𿆅6XsdF~��aQ���"q�ߏL����d�5����`K*��I�c�Z��"q�ߺ!`�u�!jJHn��z��nw=�����7`����"q��gD�+��I��'��L�m�M��T�J�Z;5B5Y+��))��wɋ��ă�s0�7��65�������uo����}��5����`K�$�Y��1�\3�#j<��#���������^P/��Ij b�S�^��d&3�-��_�.K>�5����`K�������߈�vJVt�l�褻�svJ����2*�JHn��z���NM�Gs�b�a�	N���a-��}g��u"��*�ΊJ�b����s`h�-���K�vV��B%���O|�3�d(]�/{��l�ʠ8�j�'n�^0oOH���NYY�Z�s�m�.��H�c��1�%�e��G�bZ�U�Eʃ�5�"�r�~G��;ؔ��r�C¦�bL!�DU}��s�'��U'j���%�a����.T>��Y!Ⅲ1D�14�~�Xo��0���$��c�����`�Wr���n�:.��R$��n�3R��jH�3�Ӻ��L�9G�I�j�[�.(+��S�*���X:�*��ܟ��/�b��ަ�"�K�b��Ub�ۙD���*
�I��'�:�u�J�/k� ��>f���c��1���8}�Ͼ'���ߌ[R)Ms	[�������5��G��
�O,#�N�MĐ�r�
���k�6P6x]G���i|Stߛ�D�G�
^)6��9��xx�rDc�5��ja~��j.o�c�\.U1+]i�V��`h�-�����!�(��~��j.o�ѱ}����S_BR���U�'���Xw�j�7��[�.(+��S�*���X:�*��ܟ�*��T�����Cҷ��enɌ�����14�~�Xom�q������ś���� 8axh�O�W
�������Y1����. H��z���8�ϑ��[�֊�Dfd�˃0�lS<orǟD�uiL${?�����>��yܛ�	��|��	(���<�:�9��19TH���'�3�$ �#^�Vn�^ֻ��!� c�"�;�4�t=�j�.�/'�����W;5B5Y+��A�DlO�
� �F�=D�[ \��ݪ�򈟔^ֻ������#�����$�R�n�9j�ʛ�q:i@_��u�Z����N-6�m~G��;ؔ��r�C©���+7}F�sDE�: k�g�x�s]���uC#����
p��#�}F�sDE�:�&8���l�mq���)�:��j8HQ��e�z���V�RDFR7������`��I�t?�_��B�e�D�*�Y�p�Yч���Ҟ�+�����P�[�&���_������������|�sd���C�"��T�KL�IO�!iU����jL�U���;�A+b��[	��[�w!� c�"�;���<����Dg��y��tq��*��|`�|R�:
��\|��eA&��9��k!�7�D�>����B�Vί��C���1&&��~�4�)L�sj|~��A�!`�u�!j�4I^J<�ƫ��t �X5a
\��a\Y����_�G��Gjݭ�F����/�J�Ǟ~���;���Ɏ�Ɉf�=K�4	G����7�X����Rm�Ƈ��ݱk4# `�}P��Nʆ�In��t,JQ������z��>x��F�\Mf���9��Y�{'%s�e�.YME�OW�fL��@%W�D�3����h������<�:�9��19TH���`]�n�p�'��-d�Ry��\�v����e1��N/����L�zl���y���ܴ�&�-6�Qkw�<��hθ�������PPV��"tXۓښ-x�]�V��k����w��V%�piS�G���w5��P���P���Pz����������-6�Qkw�<����y�]E� o��*�2>�1$��_w���<�Uq{�f��aƢ��K�Տx���1�|�c��1��o��yJ���ц��<�:�9������ݧG �ŴP��Cn���}/�x�]�V���HN���Mc�����n�=1�RR�,�*Ǚ62�4�ͻs�	Õ�)X�J"��Q����ʳ�A~�0 �i7�sp>O;3<�U�C��z����Ջ�/Cp�14�~�Xo��0���$��c����zL͊�q���19TH��ݧG �ŴP��Cn^�\���ĉq�p�F><1����"9o"qP�U� ���_~�?���vl�+��3�-�#���[���)gΔc�G���`NO}F�sDE�:�C&�����&� LK�a���1���.>/-ƚ��s���f���!��Z�-��AuFT���č�Y���S�)37J*u�v3���?B]z�����B*�2���u���d��O�Z�:����!n�������s�3�t8��5���dq��ٜ�U�n~q_3#ڸZ鎬�����r44���ڶ�|ceJ�z��eUh%>�L��ѥ�"���$v�~������]�!�����#e;7mg�o�b"�3�-�y�xUq�1T��8�ߒ&ˣb�O�P���H���g-�B'Ő�t(�ƺX�Y���[JQD<��z��}拋ġC����,5�<��s��]b_3#ڸZ鎬����+@�oS��7A�k�6�Ц�V�2K2S�)37J*uXm:v ��H����*�E��M@3%�?b���-(S�)37J*u����8d�^{����z��n��7�|��].��'���Xw_�'�����7A�k�6�Ц�V�2K2S�)37J*u'H?�׳�#8���Hm�č�Y���S�)37J*uV��4����?GQ�.��V��?ojʣ='Xhy f�Lu�ms|d_!�\�<��z��}�0z�cULY�ï��Jf`�g�W�����h�ׯ%�O
�_�Z)��ѫ���;����Ew(�A{d�F��M�9W2�R�E$OK�/�,�	��E"Z���Q�rۤG�#r,�-�_�G�x�J�<��z��}�צ:�)ݓ�4�A��Q�
_�J�g��0#��=��DψZ���d���-ݿL�)�y�H�������B �n�6ӌ�Iۏ��t>W��ҋX������S8���{>�JaU�C��z����1��t_Ma�~�Ǔ8���/�u�L�K4�u��t�&6ӌ�Iۏ8��0�u9�����`�^���}ɤ���
�?<pI$��g7�S�)37J*u�v3���?[+pg&1�����Z�^�\�V�n���3�6�M��4�	��:/�ҹSS�)37J*u�v3���?d�_C�Ve8�m����{��x�������mť�U�ZG��}0����ooF�!ݒ)2����x�yf��i��]�!����=o'Oؒ�b܉���i�kL�5N�6�vg;Je'���Xw��4L2�����c-(���X$�{�b�@IE�U��@�ڗe'7������qk�	(���[��k�7G#+��Q2�+�Y�T���+«7SŞ�Ӣ��WT�j
�I��w��,c�A�L')��7����0�7��65�&H�[&-n�g��U-�e�˃�����DΦ��t�?��1�TD���rs�i�ק)"�僁����7!^�V]��}R�wX��0/zﴚ��I\CZ]���O�k�Tu�@IE�U����S8�r�:-�����`y�����-x�~}d��p'k��o��`��[� ���]�!��	Ǹ�y85�s�s��
�#��W+Δ}M��R���^�V]��}R�wX�ձ����h=�I������P
7G#+�ǟ
��|�6|�+�� VU+I�eC��D>����S�� B<���J��<��%�����W(�,\ަ�It1�%n�@��V�����Ͱ���*U�&yy�����y�]֡�\�<7�X�e��ښ�s���I���b���%xI�ac�PƐt
����������Ψ��F�x`��:����gyE�sO�I�+��Ψ��FCF���y7N/����L�zl���y3B]\�#������]��������0�BE�9Y}��Pܴ��4]�Y0�p�)+�x���1�|�c��1�u�K|]�����yd�9�&���=���a_G�v�伢���/]��.�m[+Qd�/#~��'���Xw�+u>�F�+ž,�	v�]�!��\��g�X:���
,5�b'���XwN�U�R��7���N��'���Xw.9�	3�/���jbPh�`�ewU�'���Xwg�y�ޥ-jLa���a�G9�O��]�!���<J\�(y1�x�"7G#+�Ǘ0z�cUL�n����4��b��nw;��ߪ��w������H\WC,�Y>�R�7G#+��Q2�+�Yɪ}�)���x�h�6Q�7��51f�ڻ�]�!��	Ǹ�y85�k�۾�ɞ	:�
���O�g��U-�e^������?
�����<�%�y��Y�{'%s=ͱu��̦�"�K�b��Ub�ۙD��"X��[�`�L�i�-�5�H�^��gk��S�)37J*u)T{6T'��Q8� Lڈ�|���{l�f|�ό���.�Dk��v�A�x9�5�LU%����f��6�vg;Je'���Xw�j�7��`�|��K�z��n;sǳǦ�"�K�b��Ub�ۙD^�V]��}R�wX��)s[�3��k�G������4��X re��]�!��	Ǹ�y85�6i� :��O��['���������Y,0=]^	�&������y�J�#z���6B\�6�vg;Je'���Xw�j�7��o�${U��w�X�|0��X��������`y�����L�o�!� f�Lu�m�k]m���6�vg;Je'���Xw�j�7��o�${U��w�X�|0��X��������`y���0�wg%c��Y^8�����F��٬[�I��w��,)T{6T'�h�6Q�7�$���8tV7G#+��Q2�+�Y�0/zﴚ�:�L��?�<O�����(�
t��Y�{'%s���'����-��qs�VYp��HM�e��`y�����L�o�!�0Q���g���C1zho)��
�7G#+�Ǘ0z�cUL�n����4��b��nw;��ߪ��w������0���7�0>�Q�k^�ïw��O�$F���9�dMbZ鎬����/���B։��W�>y�۠����(k�:7\s�UI��w��,2�)�L����U�p��
���)�b���"v�IȀp/x�ݐ�����P���hڋ�v^�n��R/#٤M�i.�K�p}��dE���f׿���$	n��s�xՉ�T�Ұ>D�c�lQKݗZ:���'n�^0o����y�]֡�\�<7�X�e���V!���IÙ=�H�]ƭ��&d&(C�#�7#^�Vn�^ֻ����XP���$�)���>�;6W��y�3�Y�`�_������'�7Z��,�;#0L�����@�)N��B�)Yh3;C$�-��qs�VY���ܴ�&ч_����l���v�&E��t�)�8	�p���3Ns:r�vbF��@�����>��R>Gn�
�;5B5Y+��4"�I<a��ӳ�Y�
�U�q��&�_����F��@����T�J�Z�;ۂ���j_ R�ϸX��-��:�5Ӡ���5��8�t��\�v�w5��1�\3�#j<��#�0�����(_�<��}�#8K�\�p!|T���;ۂ���d���i#@���%&p&ĩ+�.q̈n�]g�bqJ��3���L}�q����iMԲ����!n}y���q���U�.q̈n�*�� �>����t�W_3#ڸZ鎬�������i.ׯ�n��B��X��T�٥��T�����S�(�I�y.͸|��].��'���XwZ�֢t��FC5��v�c�.[K��m��[-y��i�^��F
f�M���5^sJ�UF���B�D�U{��,�#�w{:_3#ڸZ鎬�����S�#���:uS�4q�
��n��7��!n}y���q���U��W�*�� f������s��]b�|��].��'���XwB��h?�J�7A�k�6�Ц�V�2K2S�)37J*u)T{6T'�Lq���Bl$P�ĝ���1��P�߭�ҋX����`H����С��J��^��y}$��rѮ�7]��!n}y��Y�{'%s2�ew���ӳ�Y�
�ߪ��wUg�)!eT<�6�Q=(�^�H��x� H=��B*�2����L\ ү��o�  0Y�w������R��a:߻�%�q��{l�f|��rs�i��=29��a&3�-��_�owђN�~R�wX��$��X>j����{�^�X�;٬sf.�7�Sx��~�@IE�U����S8�^�8��nG�`�|��K�z&H�[&-n�g��U-�e��!��'�����Vem.��;٬sf.�7�Sx��~�@IE�U����S8��(x��^;���>���l�Lɼ�,0=]^	�&������2��T
Ƨe7��
`����0�E>���9�dMbZ鎬����	�+9��\0/zﴚ�:�L��?�<O����!n}y��Y�{'%s�O��W��[�$��X�l�Lɼ�,0=]^	�&������>����'�r��'qm�±��m|� �_W�0�]�!��	Ǹ�y85�}�-���O��g���ޔ�h���o�8���/�����/�����XQ �Kk�2�J�Gz%�S�S�)37J*u�8$�O�LV>\��p}�	��D܂�A�ϑ��[���5�P3 C�0Q���g�/=ӾɎ�x���� �~��Z2��u�>��{=��[^T�d&(C�#�7#^�Vnq{�f��a�:&�>��sU�U�w=� ?����QJHn��z�n�w6��R�����&��>����:++�����Ur��R!I�fX�x%}��1.�@�Ȼ��M����}�K�
�4l�G�pޚY�i}%_3#ڸZ鎬�������(�����CcO^Z}��"X��[�`�L�i�GV��y�&_3#ڸZ鎬������e��9���b\��!n}y���q���U����c)0k"�Ι�y�Ң�{l�f|�ό���.�{�:���g��č�Y���S�)37J*u)T{6T'����f����|��].��'���Xw＼.o�Þ�7P��T�<��z��}�Q2�+�Y���R"@ПWT�j
�I��w��,���|HH9M\��e���S������
�Zb���GMVx���� ����:x�$�N�1z@�o	�Au�%]��g��xՉ�T�Ұ>D�c�lQKݗZ:���'n�^0o����y�]֡�\�<7�X�e���V!���IÙ=�H�]ƭ��&d&(C�#�7#^�Vn�^ֻ����XP���^xі�g��q������/ E�~ (�|��].��'���Xwbq,�nRT+���i�+'���Xw��`j���E�6�vg;Je'���Xw>\��p}�	��D܂�A�ϑ��[��)#�N���e�Z%�X�㊊i����]���'d��s�KT�����bp�܄��� M[B�����'���Xw;[��b��pw��˷���d�φ���;/��.���w��S�[�QTߨ�O3����KCgpzl��a�� �܈~\�Mf���9���q���U��OZ+L���Ļ���p�T8Oܡ�����/�/��Ө�2�ɤN���C_J�g�9��m���=+��.���'���Xw��F$
�u��}�xr��U�Kf�r��y@^ժ����������d�٣�����6>��T�����D��|$w���=Y��_Q2�+�Y�s��j�ŉ̯�l��ljT%q�#��]�!���1����m{���1H����Ig`iZ鎬����Y�V��#q
nː����[B�����'���Xwa'�<� \c��`ʗ�Mf���9���q���U�pzl��a��SF���v�Sx�lޞ�ό���.���K�Q����-/�Sx�lޞ�ό���.�ҋ�?��5��D���X�R�*��}A��寔ݾNt�Y*�wX8���R�Xe��������A�e�]�!��	Ǹ�y85�ӓ��������@	Q��"X��[�Gn�k��b}`B�̥���Z �W�x+Q�*c�G���A@^7&ģM�&yy���S��S�Ib����rs�i��=29��aS��na9�tT�~eFGz�T�\ ���|.�Tӏq�M腐64S�jئ`��l����u�Ew爫� ����Z �W�x+Q�*"�u	.Y��A+b����ʘ��"l�;�w���%�����DRŔ�rUq��ɤa��)gΔc�߼������T�\ ���Yz�Sk��m�S���_A���e���A@�r$T�]W��5rt,?���;��9/���`ދ2M�7�P�F�x�ˏ8[$0��h�Ezz�d�٣��c�A�L'�f?S�$�R�n�Wǖg3ȓ8���/�a'�<� \�/刲�Z���H~Mf���9���q���U��'�*3 ��H�.	OH�4k��"H$�DZ� C�C�.�.���s�Ո:�L��?�<O�����=Y��_�0z�cUL���a��N��_����b��nw;��ߪ��w�������)�`E5�'�r��'qm�±��m|7�7y�]���J����`Y�{'%s=ͱu��������T�-��qs�VYp��HM�e��`y���pzl��a��*���d��4D���t���}�]��]�!���1����m�KU�����1�G�Qc�I����1��?\��d�٣�����6>��rD�9���#mԃw���k]m��Sx�lޞ��rs�i�̚irZ%�����+�?��g���ޔ�owђN�~R�wX����K�Q��&���'b�'=�(_��Ym�@%Z鎬�������(������7`����"q��:�
���O�g��U-�e5��e6²�KU����L��Z�N3�L�t��nSx�lޞ��rs�i�̚irZ%���㳧ٍg��X����o����;e5V�]CSK�p��jO�����\�a(􆿳���Qs����b02�OtO��F'ot#�r��8��Q3U�eT(Y�{'%s=ͱu���TJ�ov� :�
���O�g��U-�e5��e6²�!`����0Q���g���C1zho)��
�Z鎬�������(�����"��a\Y����t_-Z��T�\ ���|.�Tӏ�'_@a���1�G�Qc�k]m����=Y��_�0z�cUL���a��N��_����b��nw;��ߪ��w������u��Y'G�v|�ˑ����p|3�JR����]�!���1����m�KU����L��Z�N3MF��7��ﻋ-���C�M��N��+w�7���\(FK�4�XQ Z�Sx�lޞ�ό���.ӮF��
o�����ap���Z�-��ݾNt�Y</x/��(�T���M0��1_$	mZ鎬�������(���R2�sW��t_-Z��T�\ ���D�YO���3`��s#A�w �Ǝ͂a�Z���_�q5�ˉ��@��U�b!�FwvN�S���!#�[#����W]��B�_�+�)��� Y�b��]�ٻ�q���U��,���ΞF-�+I�Ygb��dN����B���pzl��a�9g�M�G�nE�̜��W�J�!�Ӑ���<xmZ鎬�����"I����7� ;�o�;���1�忺�4`U�j�"i��rM�+$OF>�X�"�I_$\�j�V��vXę����'���Xw<��Ò\ŦP41�b����х����%�8Rڽ���b��Ո�Q�6����{M�ࠐﻋ-����2�77�E7.N�ӃH��f���][����A���l_�t������yӀ�� $}�/�J���|w:J�d�٣���9�����Og����n��g�-��%��/A$TGQ١Ӿ�$���	kSv=ݓ��E���?��9)�
rQa�����D����'���Xwd�n]Nَ+vW.䴥�`B�)續\����'ò�������?��Q�&{��8�a�;"��PÛ�U.��͝z�C���)}���/��>Y�B�^"N���<��������'���Xw�C��b7 @ߖ�J������X%��:����l����G���?��9){�����c3�Jp����&��l]mgFĝ��Mf���9���q���U��E&l�z݉2Bͧ����{���Ah�9p,�Fr�d%��"φU��ód�Xn>��[B�����'���Xw	zSW�QO˦R.a�X1aAW4?_}���Ɔ&"�ī5�*e���*!��Uk�e~���G��[�֔/$D�[4-������D����R�AZ鎬����#7�*@��
�|���^�ݛ��5���"i��rM�<��zU���BD|�	Sx�lޞ��rs�i�K��.�)�1��bMI������[�Fc�k��`y���Ў������Qkgw��.:� tN����[*$���}ӗ�=����_K�RPk�`�?��<%��짐f�-���	������bpl$P�ĝ���� ��M�d�٣�����6>�����>u~d���'��bw����$�Z鎬����Y�V��#q��_�ϼ=S����oMf���9���q���U�pzl��a�ŔB�w3��s��]bSx�lޞ�ό���.���K�Q�t���(�x����oMf���9���q���U�pzl��a����������ɰ7L��]�!���1����mctN�`Gt_����o[B�����'���Xwa'�<� \�]VI��Z7A�k�6��
�]�$��'���Xwa'�<� \���q�C��n�{5��1_$	mZ鎬�������(����&�c�Sƚ�f�a(􆿳�=���Jt�@��Yxx���7�_�<T�4���v�I_E�+kg�s��]b��=Y��_��ġC��ן�@$˺/t��꫕qŧo��K�O��C�V��w:�$o��$�3V ^�
�	m���N����B��zϘ��H4�>�����A�IECN�aFG5�
N�֌Q���L5ӥ���-���f����Oo;�4�V	j��hIڊ389�E�EYZ/�2w�+��&�s�-����d��6,'�j�Qs��!��VF�;v���R�Y���?����9����w����Ք�ƞ�.���4d+/-�C�~��������5��{���r�hs��\w=��C�L�j�e��q=���{���r�hs��\w=��C�L����OS����{���r�hs��\w=��C�L�:I�\)�
��{���r�hs��\w=��C�L�K�K� &h�Qf�h3Z6&�<�
e���4述B���]zo}'�o�e�N��V���Tz(�,�lq�X�~X��*$��]`��ض7f�ï;�2B��y,��6��ƙ>����3)#��$��{� =G���;S���s򶙧�C�X]on�ǚ��d�٣�����6>��zK��i�� La���R�l�>D�d�٣�����6>���3e���;�/���jbPhrK�@<,уZ鎬����Y�V��#qhbiT�F��C�(��EZ �:���Q�ﻋ-���C�M��N�۷��;��\o!f�	�Ĳb�M� �{�ﻋ-�����S8��$�DB��Ho�${U��w�X�|0���ߪ��w������ݓ��E�� �߳G!�a�`��}��d�٣��c�A�L'؄�f�?�b�% ����ߪ��w������ݓ��E�]���>�?
�������[p$�*��ﻋ-�����S8��$�DB��Ho�${U��w�X�|0���ߪ��w�����褬Q�Uu�2�>d�ܡ�0t��ʓ�!&%�ӄOi����h2��6_�-N�@�I���a(􆿳��ȡp��'���Xwd�n]Nق�o�F�\���e�Q�mƿ�Lg�g��U-�e5��e6²��R�A0^L����X� fn�R�k�ew���m�Q|�P��r��Ήo2�>d�ܡ�0t��ʓ��� j�}*X�Ɋ�m�;Ź��'�?�j}�ﻋ-�����S8��$�DB��H�e�X�+� �{�c�vI�ߪ��w������ݓ��E�� �߳G!#I6�q�3)�_���ݢ��d�٣��c�A�L'�}�4?k�a��0�BE�9Y}��P���"X��[�z�C���*X�Ɋ�p�����4�k����d�٣��c�A�L'؄�f�?즵"�K�b��Ub�ۙD��"X��[�z�C���*X�Ɋ�p�������{j<# �� *��Z鎬�������(����o�F�\���e�Q�mƿ�Lg�g��U-�e5��e6²�!`���� f�Lu�m�k]m��Sx�lޞ��rs�i�̚irZ%��/�rŗ���zl���yp��HM�e��`y���pzl��a�˛AHCO�i�?��kR�K=s�(:G��?�U��Z鎬�������(����o�F�\���e�Q�mƿ�Lg�g��U-�e5��e6²T�bj�V�c�Y^8�����V������]�!���1����mT�bj�V�c�Y^8����ZF�V�x�!d�}�2��'���Xwa'�<� \[	sqX��I[�Gv��FSx�lޞ�ό���.���K�Q�h�6Q�7��ob!*��2}���]�!���1����mZ�M�R���'�r��'q#�� �[N0��<���Q�q���U�pzl��a�;w>`�2ݧ�&����<�U(���d�٣�����6>��b02�Og���rB[B�����'���Xw�j�7���L�m�M����7�Xk�a(􆿳���Qs��������W]��B�_�+�)���]Iΐﻋ-���C�M��N�ۭ��_zx���ɋ���C������ft��o=��]�!��	Ǹ�y85�'���[v��`�"�X���!y(~,�a(􆿳���Qs����h�k/���J��w BM��ɋ���C������ft��o=��]�!��	Ǹ�y85�'���[v��`�"�X���!y(~,�a(􆿳���Qs����rD�9����ǆ8�ҁ���A�s<�ﻋ-���C�M��N��+w�7�k��(����*k�"=��]�!��	Ǹ�y85�&&��hO[�;���_�#:�N��u������ٕ��EW�maH.E6��P�������*	+�J�e�X�+� �{�c�vI�ߪ��w������5�e`��9�=4���~;{����Sx�lޞ�ό���.���K�Qe��)��Q��:'�T�+X�U'6^Z鎬����Y�V��#qˢ���[6}MC}5

�]�$��'���Xwa'�<� \�./^H20�Cs���ﻋ-�����S8���o�tyr�fpx��p��HM�e��`y���|��{>���'_@a����ߺ2��61Y5���;�]�!���1����mB�8r\V����p^���bFg�`P	��=Y��_Q2�+�Y��׎o�|��։�s/���N��+�ﻋ-���C�M��N���%�6l���J�g����ﻋ-���C�M��N�ۥ�`V�n��gq�'���a�ʊ���=Y��_Q2�+�Y�ݓ��E����o��W�j��6$>q��tm�Կ��]�!��	Ǹ�y85�&&��hO[�;���_�#:�N��u��=��?��^�V]��}R�wX����K�Q�B �n�6ӌ�Iۏ'�TI�A��=Y��_@D���uL�3���uZ����Sh���aSmMggE��{i�et_6�>K�fV?*��4!�wM-X����6����AZ鎬�������(����mA��֜c��x�)6��9��xx�rDc��/�;���N���7a(􆿳���Qs�����P{��
��&$�^���}��Y!��]�!���1����m��o�,��ns`&Ѡ _;��i�1Sx�lޞ�ό���.Ӈ��uj�*Hq�o�d@-[�v:v�o���+���5���L����;j����>^���o���KEd��]^X0��
x-	���'�$HgL��)�J����f5i�A��I`��=J'����r
���I}}3M�C,����|#^�Vn����o[���=^��>D�c�lQ�����+�7끍J�[T�)��
�6���.�֌���<�a)�m�d�so�}a�C�ub;�;�濖n�P���g��XQ��k8�5�>�yKYQs��[�|�F��ˮ�pd�Zз���\��6�R�X�?�I��H���Kn�ǈ�s	\jb01
�;��S��y9Ez��}��H֞��� �z��w�����4L"炡t�8j�t�Y�Ij���0E���FZ���;D8���:��M�S�ᳰ��X�z���t���Xo޲G�����$7x�c >��}f]���]�w9"x�g�Hz���!Z�>��P$��j�f��>0M�<k�lw�i}4���0�H^�wr�y[�qj�15���{v��_G.B���uOܟB8�A��jeN�V�������1d��3+'P2ӡ��,����|#^�Vn�B��מ�\P�O����X�e��rl���1)�*C�8���EBy��J�z�3fGt_�z�febÆ����9.�Ύ8�qXF�����z�1�b$E�D_��Gɋ|5���F��S�?\�ڏ �6n�N�G��s!�y�������	4T���\�nƨP�ʱ:��ԝ�XLVt����G��5�&��p���P�#�|�B�X�g�i0\��.�gIt�!�����o����x�ҡ-�ّ�^ $� 'fa�#�i~0!�r�qU���Qv�EoO�؁'/B{�;4fx��V$�w�}MX�]y�y�3�˝��28Zlۨ�\�"ߗt$��6�iy��7I��XG��]�w9"x�g�Hz���MN����!I/�������A��1��+�W�Ń�I��-NdRg�/�mC ۸���9��;9k#:̧�	��U;.��=IN�ƫѦ��2�����Vc2�����VcIv��,7�x�n	������EK�N�1�� ��2�����Vc�cRq>h���=��� ��WHBפc2���5u�OEֶ�"�b��V��;� �µ

��0��᭖K��"h��3c/��!���z{J�۞h�G�lF�ĸJ�<�&0H�N���6
�8a�w�C>��K{�R�$�V֌#V��u9z#��8h� t�э�]�,c��k�-�����qN��f��6&1�� B+@��i�s��GF�DZܤ�j<�`�hE�RǷe�b��1j�L�uVBv[2�j�f�;�>)ʐ|5Uκ��r��`���e�H�j��y��H�W۞h�G�
�蛺��r��`���9$��\��h7�a��c�,�[`�Qb��~���y���������DZܤ�j<�`�hE�c,W� K91j�L�uVB��=��|S���I�&�`��\��K��A!�?2���L�b3N��wm��5�;�H���oՖ�zA!�?2���L�b3N�B�����f�;�>)�� �4"���B�V�:��Ԕr!��I\+�U��~mVx�'�8S�E�����5�2D�3����hY���v`?�d���&�I`o����"�I_$\���`���O�s�)];I�!��I\+��o���9B<0�����|�+��?�d���&��9��^K��c��>���|�P(��25� �$�J���7�����{^����|�%����0�3p,��ùd���M���Z���BT
E7�Ո�Q�6칖�2�m�5�a�M7���Ո�Q�6�yP��C��?�;�\�R/;��|B������d���,�rK.�`�dy�V�{��\|��Ea+a�G3�u]˴�����x��ֹըQ��kGQ��l�4��H��[)�ٽ�f퀔������	-$ߔ���e�cN�V�\���vM�m�rl5v�I�D���t�:��ȝG�]��#D\�qF��%��ό�;�LȫԷ�/�P,&�ͦ���X0�6�4q̆8: D�4P���7ܬX�"������r���aM"�������M=�`�㚽6���Ӻ��L�~�y�ю�?z�:Y����*���Э��v���v���ԿK�^V�$\�6Þ��V��;��|B�`E]4��0r(�ݏ���k�	�dĭhO�^u!뼤Ÿg8V#��4�x&ʕ#;���{^���B%���O-�#���[�t
ZZKݕ�a�]�M��̋8��s�kGQ��l�4��H���0�0�h��#g�k��`�
}:�������]��:s+���6{�ZV��	��y�r��(V%����]��$^ t�ٱ"::i�(�\Dˉ���N���7��>�2�@���������B���eJ�7����K��D�e|�L�:�;�T���d�����)k��?(�Q�M�X�j�9�I����jcҦo7A�k�6��9R�$P|g��D��l��z�͉"_� N��r*\=�~ o8�1�R�*���M�,������3~I/��\]N��<Ri*�SG@ 7A�k�6����xtF�!���Fi����o�`��	����f��M�n�cqgF/�}q���V�2�C�Wz���_�%�y�%�э�����$57O��4'��7�OT�,��5�"�r�~G��;ؔ��r�C���$�&V�B%���O|�3�d(]�/{��l�ƶ�~b�!jS&�7G�hM��{ ��Ʋ��1O���ełG֨˜��C��f��M�n�cqgF=��PE���(�V�ܼ���s���LFC7�5$�)�vx�+]��ٶ����x�F�"�������d���X�����K[ҩ:�y��$�R�n,�	�X��Ɠs���^C��7cd	ACDCx��-��߂��g�K�
�湅���;��Ry�*v�FdG@9��<�l�gFĝ��x��-�/��γ�{�����F r��)�S�t��d[E�������is[�EV@Hb^�G��l=Э��َm�.��H�c��1�u�K|]����J�nt�UY=��ͥUAV�?���?��9)����`\F���%;�L��?��9)�
rQa���Hu����i&�L4⭦�����.ƶ�~b�!j�m�.��H�$��=��$�R�nl�;�w���PͿaMD`�o��>P��U2�J�D�;&Q0��6j�"Hs�VV�a|�E�j���PU�>���l�E���M��� �w�h�7ܬX�"���"�K�b=�Z��}����ޙ��] ,?I-�ǎ؎B�����r���aM"���������u���?�d���&�nPk���dDz?��\TL��E�]&I�#�P��Ʋ��1OVz�v@��'qi�á[�6���l �����4���ʽ�n8`ݧG �Ŵ
"4F��l���D��q&��k�S�|�+��?�d���&��e�/�,�g8V#��4�S��@z��אԣ#Caa��%3�xw���A�d�x� �q0)g�:jA_���t��j�j����t� VU+I��5�6���e�cNơ�&Y��V� o������ �w���z�}��g0�!�'��X�����Y��g�0�uY!+����j�Ï��	��B� �v1r��_.�yE"�B���zc`o�E��sY:�;S~�����o۪	�}a�]�w%�oφ��<�6���;�7*'��h�\w��;�jz�(�Z��8dhY�#���n���X(��;��~9,�1�12�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��Y7�0�(#;�b�`� ��I��`�S-$m��m��b�?ޓ㫝��LB�S����8]�Qŀt2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��)��o�w/D�Ù
���e?d\�2ݠ�qSJ�k��7�փ�G�#�j4Or�����g�0�u�8�ߧ\����W �-g	�X��d��S�!g�d��������\����A@�݄���Zj���������e85��_ۑ;�.IDF��eJ���i�[Y5̹���Z8!n��F��5ߧE4��Fi��|�3;c�<j��kef��?a��?cܝ\�C E���{^���l�4��H���ւ���z�����Ш;��|B* ^���x�j�9�I��&,Ξ._�0h�5e��8�ߧ\����W �-g	�X��d��S�!g�d�!��(��M�5t��v�݄�������
�?<$*K���z׏�����MFi��|ր���5V��	��yO8S��%�ѥ����R�9zY�hd�ً�e���$���{^���l�4��H���ւ���z�,�#�*z�;��|B��R����.IDF��e��mˊ��ՙ�xsq��?�d���&�0���v`�2�����Vc2�����Vc�cRq>h���`ȉ�d�M���5^s%�4�m�@:� 3l*��2�����Vc2�����Vc2�����Vc?��Q�(�'�Hm��1�dR�L��G�<p���|'�'���e�)�*C�8؉b�'��(�~��e�.5�����OI�.�������G�+Jg���]
!n)����w&#7���ʫ;�R�I͗�'7��?a�Lc�TH������7��ia1�g��M���5^s���0��_���誸|v�Q�$�W=<����c����`y����#c8o7C?����o/!�f�u�!P���b6�T��ԕ�]!B���j>��?&��Sa�4o�̽�o��`|�9�)h�A�p���|��,���ڋC�#�˛m#%��짐�CY
-����hB?�F|E�X�j:%�8� Yd���'��b� o���YdZ0o�v��?B����ߍ����Nu���[�9]�ܔ��f�����o/!�f�u�!P���b6�T��ԕ�]!B���jc�|M;�~M�C:4��7A�k�6���u�iX$�M���5^s�F�O^1�e�^#�6����Q��\��k�"�RF]7A�k�6���u�iX$�M���5^s�F�O^1�e�^#�6����.B�M޺��Og?6������o/!�f�u�!P���b6�T��ԕ�]!B���j���7����KP�	��k�!!ʽ; ��#f(Y��[�n�{5�aX��;�x��B#ݧ{0O�}����h(����F�!���Fi����ot�*hH����.^݂�`� �(��2,�<I�Cl�6j�V��vݟ=�NM�zk�����7�Ѵ���I�q(��h��4NV�e��1������Ӻ��L�~�y�ю�?z�:Y���IBN!�e�[(7lփ�G�#�j����u���SYuN�Ū|u�?b�L���dL7A�k�6��K��8{��b�&�q��ax��Y�L%�z�-uͺI�s�U�q���5X��WG ��k\R�g��:��T��ccd`�.ۗ�臣�4}���9H�f	$��gU-���
G�|�!<��/�ciJ��V���i_r�(�������b�������*�
�ؗ����$�j��:=�����tg?_��{�f�d���'��b��oS���*�M8Z�,�\�)�`"���b���f���fa��[��q{mB!�����ɣ#�fp�J��{A����a-6�Da!��I\+��o���9B<0�����'�^����#k�˟ܒ�o|k�Lb�5ߧE4��\�ܢ��,	սL��$����,�ǰ�!@� ��Z�b�8�rW6|Ǚ���v�3�&��p�E"�%|9�1	��e��Żl5v�I�D���t�:��Zcqe�+�;��|B��W��$~�I`o����"�I_$\�j�V��vݟ=�NM��IC�oH��;��|B]it7O����m�s�_�~�)#2�����Vc2�����Vc2�����Vc��Y7�.C��6��sNb�ۄ+�lX҉N8*֑���2�����Vc2�����Vc2�����Vc��G�ZB���cp:��G�`��K������� ���9#�35xM�����?��9)HU�g���nF�o�F�w����?��;�Ӏׅ�S6Q�8��A���-s��*3M��t�[��(�2����0�s��# 툻��z�~�����8OT��)Ø�O�qPl�W˝�ѷ%��짐"nq���z��Ӯ��N����5F��U�B!'ћ�}��`�K���=���o�8[k؊IP�����hJ� ��ׁ�R�o{�}�`��1����;� v�ȧ�b�	C�d�&j�>�$2�N�9`�p�0|��0����mp��{ܤ��A�g�/H�|N�w?���p̦/�:to��h�T��*^�8�k˄�K���zռA���K�MvM�u��8*t r�D}�C7F�=j�=��Ѐ�Sn�d����6�_z��������0��&T�ͪ͌�>��Tz�	����i�b��3K�<�BJ�gwr���iț�1?�>���^�����K��^�.@ ������e �ǟ=EZF��S�(57^�	���ry�TG��~��]^!�U�����CͲ����9h�A�t�+_�dG�y#�
A�e�:���D=,Ϩ4���� 	�oݦ��D��ܒ���JlwL��{��L�ME�E����>ˌ#�0ۙ���-!^�����K�����i{��W��(����ѕ��J��<�..�4��\��������ώM:��2�,����|#^�Vn�����'MB�I:׷�Fy�XZ@po��*���3m��U}�	�2�G�Ml\P�O����X�e���&qL�+.�/'�����WX�*�܁�c�PƐt
y�XZ@poI�H/�v�6���l �?��CGqi�á[�6���l �M���&�=D�[ \��ݪ�򈟈�f��2R�A+b����)�yI�H/�vŤl��%�_���	��f�[<��Md�x�s]���uC#���:pw05TS��t��)�����)9�[ƅ���H�VF-|��S��t��)�����)9�cel��oW�7γҬ�,;���ʘ��"l�;�w���\���L>�l�4��H���F(�E����.�x�� E^����<b  �H�,3�V���C�m��
���)^>�b*b  �H�,3�V���C�7
W��;��Tɀ��T�J�Z��K�Ō1T��v�ܾ�y�j\��QםJ e�g���ޔ���SS����F�xE�W`�|��K�z�)�p*��L�+�M�R��x���hÁ	P6���N�h���.��f�M�ވ�'��Ǵ�X�)Х��㵾�Fz� �ZBh�Y!Ⅲ1D�14�~�Xo��0���l�2q;H�-ވ�'��Ǵϴ`�-2c��ҭ��'���ߌ[��83�$^й��Qm�N�߄�4�X�)Х���[� Ag��g��U-�e[�.(+��S�*���X:�*��ܟ�� J�&/��>�SS�]��Rm�Ƈ��ݱk4# X���|6�k�#��.���t�:�6[��j��(t�	��i|Stߛ��ȉ26���\P�/vփZ���0�́	P6����`]�n�p��#��rܦ�"�K�b��Ub�ۙD��f��2R/�rŗ���zl���y��(����4&ݞ9����F�4B�[ƅ���H��*�5�ٻ��E9k��-��g<�*-�RԚf�4&ݞ9��h�xm��.�3���l��́	P6����4&ݞ9��h�xm��.�3���l��5��U�߈�vJVt�l�褻�sv�J��
�D��j��'���MIM�աRC U�<��zɛ����|�bІ��xx�rDc�O��Юlb�1���v�)6��9��xx�rDc�ቩW<$�X�~*�R��1�RR�,�*Ǚ62嫐��r(�X��+�p�U�C��z����7��j�5��½ɋYiݧG �ŴP��Cnլ���4�L�U���;��n�^-p��G-��\)6��9��xx�rDc�;��k�Q�C�������P'Q^�(�]�*�|�bІ��xx�rDc�E|s���J���l���8��!����eQ?��*�5�ٻ1�RR�,�*Ǚ62�y��{W(3���P�5��$�/-�!��bk1�RR�,�*Ǚ62嫫�Rm�Ƈ��ݱk4# ��sw�r��8H���b���&<U�C��z����Ջ�/Cp�14�~�Xo��0���l�2q;H�-vl�+��3�-�#���[���)gΔc�oG���g�)6��9��xx�rDc�虎لN*c�p��I���p&Zc��gc�jv�Тk���aA�h�Ӆ��x��_���wg�W���'h���W^������h4c�Ү@;���!ѥ�"���$��v·��.��6�S������R]Yp���Vh?�����=!�Ca!T_07l�"b��"am��%�t�B=4�����o2�:�r�7A�k�6����&�nP{Vf����aUZ���RT�0]���!Vf����aU�a����:��$�n�-'�(�����Q�_�N�g�w�����7A�k�6����&�nP{T���M0�E���Xyܽ�޹ܮ�W7A�k�6����&�nP{s@�&eVC�����+H�K��J<W�f�ӊ[�k�T�"2o����\�o-�Qd�|��aK ~ж� ��%����
�?<�K���SN�b'&�3hǴ�� #��L��_�wb�md�����H~ �
4 �g[[%씡��j�ӂsZe=�|�:c�]Dz?��\T\Y��ä �m�@�?FZ�±��m�^p+�b��Z�������u��w1j���!L#�]2 �m�@�?FZ�±��m>˟N�0D-��K�}i�R���O�C;=B>�)3����ՀW�l�l���XU(�a�0/zﴚ�/����h#�88y�[��e�|��ooF�!ݒ)2����x�s�a�p梯�DΦ��tL��,c3ಙ��%!�t����V���0�wg%c�_j��r�.%�H��,��YzoM�B8�\�W�EC����pLC���� �%�H��,ۙ��*Ը�y["�W��@`EE��o8��������)��[6�����H��:Y3Iz�SŞ�Ӣ��W�7~J�>�h$G�����=���+Hx�/�l?
�A���g�8&f#��։�s/�? �t�a���;V�����
�?<l
b���M��nq�p>W< |�;�Ojz�Qr�{S�$�:���N3!�U\���<��
��P�m�С��J��?4���R;� �U1]	���`Zf�Q�@��߿c�!;�a��/8���Q>�^2�����Vc2�����Vcv�iL�D�6,��K�d�Q�7)�G!@)c���Fu)n2�����Vc2�����Vc2�����Vc���@�	�,G��tn�U��o�������*TK���[T� t���|ӊ�.A�_�y��Ld_ ��,*\IJZ�f�$�C���J����Usr�u}��Y�&i�b�
úy��Ld_
.�Ʌꘔ��jH�X��SP9�=������i1��s�$�����)#���d/Z ��P��$78�ڠ!��2�[�'e���ܑ�J��fW��n���#B�׺�s�B��%��"�󇦕T��6ܭ�e��:s*�&*�K��|Y= D��ma9���$H�[<���9��̵��C3�']@q�5dV��$V�k��	b��F�s�����zFCHc�Me׸��R���pG/@_8�
���9*�E1���e�P���x�&aZ�+%���m�&�_�E����ݜ/�"E�m7_�ѷ�m{�HCڰ����	��D9s{��OQGT��v�F#�5�����c�_v�F8o)���,�3O%�g��!Rf��͕��:�.��ճ;$t��9&:�֖�֯��q�Z�ȕ����LT��B��7��@,�hn$�E�#s�8FTy��0q�\���wu�B*�2������Ȃ�(��F��[�}��&v.ho�Bĥݜhu��$�?8q�ש��/�Pc��?@W��7�65��{�s�j��۽b��PCb"׏+5'��Y�U�fGm��^�J�w&��)�δ�P�-�H/t�:��8C��gK���V�<R��5��!�ǟ:��'�5kPc��?@W�����9��)�A� v��F*c����bؗש��/��Hti·/7�'\�"��󗼶M
@�ͰY�����P�|S)a�q�|�O{N�M�b9��-N��&dF�D.�1o���{3t�6�2~9��g���hu�`�6d.��HP[�$�����g���?���CL�
�7�Q������\�"ߗt��E �_�N��e��!s�x��X����6�O�jB�ݔ�]<��	(�H�QbY^F <=ޮ�Y��Nv�q_X��ղ�J�)]�O�_r �:ys!�Ǐ�n9�t��B$~VM�@i�����	����(�{xt�4Z�U�W�����PC�ZE(_�>.����w�?��?h�l8QX����}0x�yZM����5�Y�w����Țuٳd?��B 䤛;m������F����x	ԛ���9������ B�h2��=-sЗ�x�����诌Q)�R]\�Y��w{��Z�x>x�0�(�D��U *�f�}ݜtR�.ǻ�rx'G���_����^lc�.[K��m᳤��5K/���	B�]w�Rd�����!f$��s�By}Vːs=3]@ޞ�޳��k�`���D�$l�TE����o���̫5�Y�w����~W�����6�O�j{�u����9��F��6�-�|��2"c�pJ^l'�J<!�i�&���QP1d; k��Dr��Q
��?���:(�C)�F��-U�ɓ�i#����7S��Ro8А��By�_"� P1��r�c[T\t�z����C�j�����ፕBH.� ��)��]g�tҬkb�H�_���a|R9�4�3���T�JdW����vJD��@�s���̴�hS}����k�l��U�X$���m��eF�m�v�R]L�Mֻ���8w�Yi.�!h����
!�]VI��Z���2M~8�#���	�}���O���'T���+��cd�1o���]�U���L�o����\�W�ECCᏼ�����w_>����	O][աI�2�y���(�1�sx�\��F����F&s;&���2nv���;��z��g�o30�A�zc��#�uRmu�/��@��0�H5MT!�J���x�z�ŏ54؋�U�a�t�o�B�7�P@��:J~�)�δ��ʘ���r}�Wq����^.�A�ڥW�`�* �*Cǁ�l�����˺�ʘ�p���ʘ���r}�Wq��*C�5(y��Y�RK����r�t\oG �O?i��{��Ǭ�s ��5��<w�-p����0<���Z�>)��	s%F'&3�˩�Ϊ���*��O�t��yoZ�P/^TA`��CSH�9��-Mq�QB���_��!���f(�@+��������\��jT�):1�#���M�zR�D�^��! k;�Pa�g"�W��{��Mm�9��� �}�; Q_� �Ezv�*J�|�U �l�2�&�^C����r��6*1���jHM�����[�g?	��o�ax��Y�L�j��SdZ4�!��Tӧ~�Q6vmI/5(Q�g�+%f���atr���pu��S�a	J/�ʵC<����P�l!AJ��w�����L�Y&D!�d���L�o�!� f�Lu�m�k]m����5�ź��\[��� f�Lu�m�k]m��g�y�ޥ-ju�u[�z����?b�%]n9��h�6Q�7������bo13�3��ŧ���X� �]v4f�D��ܳ�J� �߳G!�ȅ
��5u�>����9��0Y d��M'�F2���}���ݼ��1�G�Qc�`_���pRW�!�
�ڤ�1�G�Qc�I���З������;��W�& :�L������d�С��J��:�L���v1a{J��������;��W�& :�L��MN*����h�x#�L_�(D{ͬ�y�4����H|r��2�����Vc2�����Vc2�����Vc2�����VcIv��,7�x�0v{K��k��T[�x�(�䏓O(�e�C�$2�����Vc2�����Vc2�����Vc2�����Vc��3��kD\Ӭ��SG�d�����cab��f�k�8�4��Q>�q��w����,��>�[C&����*�E��M@3%����J �1x�it�ax��Y�L��x:A4bI�s�U�q �~k�%��x{^4��*m/�M۴� �Vf����aU�#�fp�J�!F�R��Lq���Bl$P�ĝ���Pع���;Ȼs���E8��5�:�^�h5���٩�Y�L,�p)�i/j���p^���Fh��'GXx(�i��/Rh�x#�L_�(D{ͬ�y�4����e����)�Շ^��j����
�?<�aYR�B�d�O�'@i��E9k�v��=ݏ�2tP���Q���FO�[�]���4�磕����
�?<l
b����r�\r/���jbPh�W�wx��k=�Cnpă�3�c���51[��wEGͶ0h�5e��8�ߧ\����W �-g	�X��d��S�!g�d���z��R��ؗ����$�j��:=#o�]�ʄǏ�h9x���yoZ�P/�����Ut�\�cI��S}HB��L�Ř>���q��ߺ2��t��A�ʛ��pP��Mb"�*�d�����caM�%�����t�'%����p^���~����r#k�˟ܒ�o|k�Lb�5ߧE4��\�ܢ��,	սL��$����,�ǰ8,�	��Jz9���5E f�Lu�m�o�u��*c%���i|7r��@�����5H�'�8S�E<�k{���� �g^M�va,�X����_�4n�c?�d���&�D�;E���q���:�!���p^����y�Բf�9g�M�G�n f�Lu�m.w[vB�0�&O�;u��M��7{��(:/�b�&�q��ax��Y�L��x:A4bI�s�U�q �~k�%��x{^4��*m�D�$0��X$�����gtv(�Va�ir�h�6Q�7���yoZ�P/�����Ut�\�cI��S}HB��L�Ř>���q��ߺ2��t��A�ʛ��pP��Mb"�*�d�����caM�%�����t�'%����p^���~����r#k�˟ܒ�o|k�Lb�5ߧE4��\�ܢ��,	սL��$����,�ǰR{~g�O"Z�#��������
�?<`��Đ1d��։�s/�e�*[�9��d�����ca�C�U2�����Vc2�����Vc2�����Vc��;����KW�*�	S,�d;vt����g: k��2�����Vc2�����Vc͞����C��m֐������e�  �.4^�&��t&��j�қjI�"��)�l�+4�]ed��{�b�IȀp/x��,Q��	}QorǟD�ui9�f?Y�OV�W|�B�I:׷�F׫�J��l� �[��׍��������֡�\�<7�X�e����]��m�n������"���P�`m��';��?2^�9<o�nïi��n�5�F�^hq��:�����Lh�7�Qa�_�G��Ǵ	P6����|��{�r�\	��rR���k�V�\���e�Q8-�^\́	P6���o�${U��w�X�|0��ѓ�s���O��['���x��U8��\���L>����e�� ������#��r������r���aM"����E֤�*�5�ٻ1�RR�,�*Ǚ62�3�����g�m>�`^����S,د�p�L������� ���8�%e��ڡ7oA!�䀯�8{+��
uj�����O�D}�����ņ�a�t��A0n���J��x��uqq9/�)�ԙ�.������Xuε�!>��/�����j"^�����ϖ [@wP=�	�:˳0ʓY+���_D�Q�C���� �
±2��h�6Q�7�0ʓY+��g�$��b܉����]I�9�\5">�E �9���=���˵k�^�pfn�R�k�ew���m�Z��-&�-�5�H�^�i�ӎL*$c�\�^>ZObW�!�
����
kX��!��ೣd5�͐��%�v�x�zIb�E�0W�l�l���XU(�a�+93��CxO�`
�-��d5�͐�-��;���:�n:G�j�jz+ ^,e(}�S�����4�֧��L_Q�����f;��V��m�;Ź��'�?�j}�˵k�^�p����X� �Sy�A-,�:���N3!�J5^�ұ�|��d��w��L9�ۘ��ҧ�?�\���3cx���K*Fg��,��˛AHCO�i�?��kR�KB��}�)�<��D�V�}Q4XʰS'F��-�x�h�6Q�7��m0n��,�0�wg%c�ִ��#"�w�Xb<���h�6Q�7�2�����0/zﴚ�:�L��?�<O���e�|���Dsw��J�����:��!$��;�s�*�:�L��?�<O�����+�	����X��֑xGVָ]���=A�%&^�nƒg�|R��qMw�}g��ti4c�St��'�r��'q#�� �[N0N�b� 0e[O��ɔ�<5���3g6�9
��G���1j|g[Ҡ(Y�u�/r��#�<���=��s��Q>�^2�����Vc2�����Vc�Z3߯���oL��ɭ�����Ni���2�2�����Vc2�����Vc�cRq>h�a�{K���6B\n���Ϩ���]k�kIY��oBd?\$��M��ݺ|��W�����ώM:��2�n�ڤ���[U�&�nЮ��\�]\���e�Q�����k�/U���!-�iP��G��\OL^��>%�Нo@���;1?�[F�9��G:([9��qUB������Wi�g���h���R���ɢ���ڠ�Q;�m��j"^�����ϖ [@wPcIn-Hzn�!��ZBV�RDFR7��D�
p���kg>�[OF�ѿa@��h���R�޶(xʶ���H3=-��7��k�VX��he�	q�X�Z-�_���mA�N�\:����v·��E;�ٺ6�w�н'�o�t��;��"h#�)��*N/�p��>E��ѸZ�����=[����ѵ�������?��ًGx�6��*B4��c	�yE�,�I��ގ	�� �\|��Ea+a�G3�u]˴�����x_��s�֙Q;��؆JWJ��w BM��ɋ���C������]��<a�9g�M�G�nE�̜��W����u�u�d!j�e{�~��j.o�ѱ}����S�U<f9^6To�${U��w�X�|0���ߪ��w�����蜗��,�ǰƺ��kÄH_��#��aѤ}[WckL(�Y��1v2��W
_F@SЙ� "̧�Y��\|��Ea+a�G3�u]+�u�G�k_��s�֙Q;��؆JWJ��w BM��ɋ���C������]��<a�9g�M�G�nE�̜��W����u�uPs_*�GqW�w��fD/����p���_V�r��%��;�tI�g?	��o���Y�]~p <�r�\���U(E�pOd<N�!�Q�f�:3b��J�Ve
�AOWm;���:Y3Iz�SŞ�Ӣ�F��������Srٌ�y��Kᷪl?
�A�� L#_/�e-M�O��~�y�J�#z�3W�ǡ¶֢��s�Kȏ���*�o!f�	�Ĳ� {�'#��T۳�͕��AKd��y c�gtb4�^���F�f�J�Z�G�O�(J��w BM��ɋ���C�����Ӌ�T"��D�x(�i��/R�������	սL��$���7'���I`����%�XDH�tt��ig}@��Q��)I��B��7c�p�V �!8�8C��z�:Y�����gڟ4���I`��y�<zQ���n��뾦��c�������C��#��>��:�@U�g�q��}.�WyT �$:�#��>��:�@U�g�B QU�Ka@��Q��)I��B��7c�p�V �pf�� i/�={"��sZ���Y�!�#��>�a$�i����c�Z�~����,�ǰ&k������ǆ8�ҁ��Tŵ�$R�i�Yl-)@xz�:e����
�?<.���6 �pN��r��<Н=.��E�E��Z�2�����Vc2�����Vc2�����Vc��Y7╙f��/(ޮT2V����uV(1тQ���3�u�l2�����Vc2�����Vc2�����Vc��`���4"�A^�F��gVE��Qx�B��������e���F�Z1��}ٲlY�T5�����=tQM�_����6��LM�<�>u��N�x��e��k�7ܬX�"�Hb^�G�𿫺}Z35�V_��s�֙C�T&L�P e�mC`���j��k{���e�V�{��$���G�"�M��.!y�O�|�5�<�..�4��\tb�Q��b�:�	$?�����e�>64[`�)6��9��xx�rDc��/�;���)�v������t^���\�}]C^�5Q��R���|�ޣ�W�]eeݐ���м{�%GuN����A@�e���?ͧ,�EXt�|p.�����4���ZU.⭾)6��9�ߺ����T�2V�q�Y�;�
��+�d��[{���_,�c$�N�1E��Zi�DЫ�5�|���XԦ,\ަ�It}�0�.�,��.0b��V�����c�,�%Dv�y �谝��X�e��}�g�{wln������Y�
� T[��m��U}�	�(��Q|3�r�^K������О.�!H6F�� .�/'�b���' /��~�;����ɝ\�!2A����ed���M��7�vsi����WG��6`Bmy;;���0��0��}���'/e����'3Ȉ�7�u��\<g�
7�����D�nR�����,�ǰN����;��Y߸I~H�1u$���B�����(�m��w��l�U�C��z��
������y��ٓA��E��锏��Z��E�ㄪ���wM-X����痴�y��������z�	q�JaQ�Hu����i&�L4⭦�����.ƶ�~b�!j�m�.��H�$��=��$�R�nl�;�w���vKz��+�c�����|�\;͖�kYIį�a�y{�הr�R_ǌ��g�0�u\=�~ o8�1�R�*���M�,������3~I/��\]��j�/A=�� ��u��ۥ<ab�۹��{q�J��pc,<v
\�W��  m�K��*`,9�H�WgＦ��Jl�4��H���F(�E���;�
��7cd	ACDCx��-��߂��g�K�
��kmٸ;͑�؈a����ry����{�Kv�]���=�n�!
����H�.�R�Xe����>S��J�"=��PE��
��T���x)W�Xo�5ߧE4��\�ܢ��,a�U�ے
�篌�	哔דo�1I6�F�,�֏�j�Ֆ5d�,\ަ�It�� �18�n�֒ce�?*h"���3�$X������㳧ٍg��X����o����;e5V�]CSK�p��jO�ٺ�oW��j\�/��Я��AS�ӡX�i��]IN��_����b��nw;�ny4�%$�J*��u���>2�ۙ�S��na9��AD��|)6��9��xx�rDc��/�;���20k��W7��c�r�"��%����$X��������+�?��g���ޔih�7�=���yp�.�-,H�
 ��X�i��]I�"�!1�U8�LC��i��E�A�r^J����'�{�IhJ�(w�Qt
�B8�1CY��;Ξ��\So-�>�6C\OL^��>%�P�^/�h�SL@�>#}��I=�=�x8@�*�p͑����5�8Cl8R�a��H�~��O�G�D���1��uO����lDx�֣F3��O�G�D���1��uO����l�^_���mo�C$���4~1��@�C,���yx�E����l���tL��4~1��0�RQ�� og�6�G�8���4����6���״��D�,��qZU'�`-�K�تG1l��)��fC��T�_/��
��Lh�7�Qa���ﴼb�<5�\��w�wF?�d�0�D�Q�~���G��cY�����Ї�J}�������EF�]�`�|��K�z��d@L�Q��d	c�b��yx�E������Ka�l��)��fC��T�_/��
��^7^�γ�4���ﴼb��|�Z`��w�2*Q=F���q�4�^7^�γ�4��12~ "�&��d��:n���+���7��
��[8{�n�_ ��n�Xw�5�8Cl8R�F݊h- g�x�&��'����;�5�8Cl8R�����E����4��Bu�(x'�2�i��F�eh���6a��bft���3y�Z0_@�C,���yx�E����l���tLC�mr�,'�0�RQ�� og�6�G�8���4��;������״��D�,�T�<D����;:\$h�ld'�V��EuX8�������=�Ҹ�S��F��u2�k���ձI���t�i��;��6�������Лz��ZϷ�@��;h���X �j0��.@.$,�ͼ��%F��5�w�|���7-]���:9&N�'�̀|�7�<t&Y_��lW�B>l�2��!�qS���T�ژ�k��\OL^��>%���Ѐ��~�;����ɝ\�!2Ak\R�g����Sܬ�T���>�M���<���2r�i)
��FP�?��ԭ�P����v�^l�}� 6ئ����3}� �[�ɦ3�pe��,!���;)��4{"(�o-��	�!��ZB�ح(��4D���t�vJ}���X�m��%c]+93��Cx&�~6�	��]8u��lm�:�L���v1a{J�4��l��������l8��P�U��<?h&�,�|SY�b�B�`zLנ�3��!��ZB�ح(���@��b�iR'�&��܏��-B��!/�H�h�c6;�L��Z�N3j$��1�#t�����l8$�LM��[�6M��Hz#mԃw��_Y�L�������l8EF��|�Ъ��=�Z���D�nR��X�ۥD!���
���c50�ś����{^�����"q���
G<�K�f>x�:	d�#��K��t%>^��VP�y����fD�b
�,%�٧�\�T����!N�~<6���Y7B�p��|(����ã��8HS̅+s���a�㑽���.�*@�� c�Q�ټ:��N�%U�0_�=2���XKa�QU�g  ��hc^�$�J	ъ)�އ��622���mg	}�î\�������S����>AU!"k�\OL^��>%�>DM��t�/s7gX���� s^r}����PATՇ�`�v��|�o�0{}i�&�a���|�csr�	ؖk�`P�	!�s�?G��TȖ����e���W�l`�݃�<��N�L�i�CͿ�����.�*@�� �]�;~�/&$��8_�/s7gX'�-%�t��y(�����������(�����;���]c0�]�:�9�sCyu,F&yh<\Bޱ�~��F���>SEL�A�;#�tױ�1�c���׭�ퟯ�Z8��f��2R�#��ٔ���y�j\�ꃤ)7��AiO觤H́	P6����e�X�+� �{�c�vIH���hVJ��|2�E�����;ym�״��D�,�w�ō���v1a{J�l`�݃�<��N�LXm�NR����0�.�*@�� ���⽀Y�k�k{����r�b�p?����z!����mg	}�î\�����>%���#g���;૞��R�[5�(��%�*ҕ/s7gX�z�KdL��h���X �Z���
�*1�3��&lk�?+aTu�z[A0q� \��l�(f���/Ax��}*���1��9�ݳ7_�Kh���R�ޭ1[�C�ߌd�r�ّM����Sq�#�-�W���G�Y�iв���N:E�W�5hG�O�] ��r{�_�ZVD�t\��s`ef�&��.�S���/�@�g�Mc��M��7�-�혉�q���z�}I��&�nP{�h�6Q�7��ob!*�1QiOͷ<e���VA��v·���Vem.��5D��0h�ky��.�"��Jg�C>���v·�<�}��O8s`ef�&���TVe:�J�2�;h��5{?�6�Xa����gB��}�)��F�D�9�lz�����|��d��`�D3���Z�/�0���/�3=M��;�YJ�� 6j�"Hs���fsK3k����O�}o{�K۬A-:���c50�ś����{^�����"q��:�CB}&��f>x�:	��)�!�B`���Vem.��5D��0h���lr�q��H��efm�0z�cUL2�H���B��j�t6j�"Hs`�0�$!�_��,�6�£p�=^���%�����jp>J@��樸Bk5G�v��&M �m�`h"�\~��MI��<2�,Dˋ�1C2,��ح(��� �����i��l�T|��c�v��N�	y�W����cW���G�����z����������ɺVE�-=�����یE�&jRl�Hm�~2��S����*�����g��ǒ,�f�*�\�c�}ڀ�V��	��y1vXD�)62�����Vc2�����Vc2�����Vcl��w&� &sG��>���>���W�b��Ǉ����Fu)n2�����Vc2�����Vc2�����Vc8m�Z�_��?��0Sߖ����Z�t���(�xx��e��k�7ܬX�"�Hb^�G�𿫺}Z35�V_��s�֙Ś����z��5�P3 C�_hAֵ��;�}C~M���p��=.,����kY��?z�٧�\�T�q�>�YŇ=�er߮�,����|#^�Vn�����'MB�I:׷�Fy�XZ@poq�_���13�[T�)���V��ÑR K�R����Uܛ�	���G�˹Ď�@���U@���:��F���Ed8���d&(C�#�7#^�VnC^���>�;6W�&[�Z�{��E��"w Wj�)��}�OV�]qr����}	�Ճ��wW�����Q:Z.�M��0�BE�nM̻�
.�2�NT��b��nw;���p���������T�-��qs�VY��2LC}��i�����y�2)����u����YcWT]�GA��"`�|��K�zSu����P$C��s���O��['���-�ｾ~:��eD�#[�f;q�s��f��2R�㳧ٍg��X����o����;e5V�]CSK�p��jO�ٺ�oWǚ���|�u�T�J�Z�?��CGTJ�ov� �:C�?p{^��D5l��i=���[&��?��
́	P6�����ӳ�Y�
����.Cih�7��fpx���:�5Ӡ������:��$�Y��1�\3�#j<��#��g.[�Tuj|~��A�!`�u�!j��  ���EW��P���VN/EI���āsp֟kh��h��#��MԲ���d��#��r0O�	>gc����h4c�&2�PK�_UE1���yh���X �a�PH�Q�t�t(�ƺX���ϓ�S	T�	��p�q�����eM�C:4��7A�k�6���MT�S�b��c�v��E���Xyܽ�'ƌF���ck�Bɉ���o��:}G6]������$s7A�k�6��G����Cl$P�ĝ�����M���̯]����↵��<��KA�E�+kg�s��]b��ORniF�!���Fi����o*��F�w*�|�1��?���HEcO�B�����{�^�X�5D��0h�ky��.�"��Og?6����@��b�O��z7��{?�6�X�R��aڊ7�C���]K�v�I��L��Z�N3?�<O�����u�Y�5#mԃw���k]m���ד�V^��\(FK��WdM4@��Z��E9�H���Vem.��;٬sf.�W�7J�Ka�t���(�x�_S1�����o�>�5�7 9>�B�5D��0h\Ef�>��t�6��B%�ɏ�X,���֑xGV�g��,��V�RDFR7�-��;���:�n:G�-}ʙLY�>0Q���g���C1zh��G���,�ӎ�Xp�,4�֧��L�q����W�7J�KaC6�=�����!���;����J��'5�S&5M�YYroE�4rh��|���W�t��m����e?�d���&�sS�"u[�T�/ֵ���=�2/���'�8S�EDy4OvvMǗbfv�\�|��Q���FDץN����v|�ˑ����p|3�l�1C��(�6{�ZV��	��y1vXD�)62�����Vc2�����Vc2�����Vcl��w&� ���@�F*>�DO(��G!@)c���Fu)n2�����Vc2�����Vc2�����Vc�Pʕ��,���Χ�0_m{��Q�'��P��+BY��9�45��\1��jHM���+t��A_���i�VJƷ7%�)�1��bMI�����5�
�J��)�1��bMI������5mݶ98��Y�d�X���l����4�n���xǊu��^���D�)��n�)�1��b��4z܂<��'Tb|�0�����&����
D�5���>��v�����&����
D�5�/�7�[��+uթ߁��N}H����	K$�ْl��]�B}Ю�0�`m��';��?2^�9<o�nïi��n�5�F�^hq��:f��3\z�[
�}3��*���1���{+%�xpp���e%(��߮�;�;�^�h�=�7��"�5h���X �Z�^6��9��tH��Ecc�,�[`�e��h��+���D�Lh���X ��f�;�>)�!�#䶜��{�:���g�h���X �4�����:�K@4I_�GZ֗~�K�ȯ���C���� 5#�3�uW���?bS�xǠ�j�!��!b��ߍ)�����߮�;����0�E>�P�'�h�&2�����Vc2�����Vc2�����Vc2�����Vc(��}�/��oM\`�)nQ �ղ2�����Vcl��w&� 2�����Vc2�����Vc2�����Vc�cRq>h��^���GB:�(��E0�gǞ����R�Q��=f׿�������!N�2��_:��y$[|�h���X �D��j��'���MIM�աRC U�<���~`�&�b�% �����s&:m�:O��['����W�
�����Tɀ�5@��>U�L�#_��,Vit�-kݔ�yN{-v\L��"��#nS#y����Y=�د�p�L�������>����V;5h���X �Z�^6�D4�ky���v·�=4���~9�n=*w��8 :��tx��az�d*�y3�/q��xZ
��+�8�K�K]9^n�Y?v�<�y3�/q���G����N��;�Ż�>%�X�Wt�MoSN�W�S/f��e�WDv�b��h�Ӆ��x�"���
wh���X �e��)�񗐔�0�E>���=��s����0+C�G���}Q4Xʰ�=�l�w[�6����'���?��7�NI>���L���dL7A�k�6��D;:dt�|:�L���½0�M����XsC�CW�[��FWv7��X>����fu!뼤Ÿg8V#��4k�z(	�����C ��X$����,�ӧ>5�L?��Vf����aU�ꚽJGrP�hG y�7㐌QjK��+�R�7@���Ӈ(j7h�4D���t���Ⱥ�����XsC�CW�[��FWv7�y���؍��9g�M�G�nʞ�sB�_\�]��"	`v~�z�xE�?F ���������l�ns`&Ѡ _;��i�1.ڒO��ikբ�{����n�bdk��������'�r��'q2I����Ċ�ъg4�֧��L_Q��������Tu�M� q��k�L'.�\&��eƀ�F��Y���j�[O��ɔ�<5���3:��m1q�cr�����ܐ�}�&��%��Bw`7��Z��u�IՏ���gN!���Lu���}Xx��(��M@3%�9tJ/.�HL���dL7A�k�6����L���h侈���&�kc�*of�����U�ӿt�xZ
��+�8�8nKQ�D�T���M0�I A6˃rG��T�J���I A6˃rG~�����0��D��l�͆��ڥ�4$��yÇ�me�g���rB��_�#��f�:3b��m1x�!z?4�e��>�\�W�EC�2[QvA�1�m�.[�}'���y�Y^8����ZF�V�x�!��*�X��j��6$>q���<��w���{^����c,�$��1�2>�1$����P�޹1�#�
_�jE^���\�}i�S�E��:c�hh��:���N3!�U\���<�y�r���,c���L�Y&�!��;�����L�Y&U%����f���5�ź�IM�P�Eݽ�"�{��,�ǰ����s�{��iK�D�b=[B� ��\ً�>��OuЙMǿI?����)�����MN�F��;���_�#:�N��u��Z���=i_��s�֙B���y3�3G���S* ��S�:�M���Cf<s0+�pΡf9��`�D3���Z�/�0��)�P؎ߤ���&�E��"+VqS?�d���&��Ln�"O��ЙMǿI?:K&�^�1����V�������t��2�����Vc2�����Vc2�����Vcl��w&� ��tF��J�����{��ܨ���[����9�GKP�2�����Vc2�����Vc2�����VcSd�*-}Q��eh��2B�k�`�?��<��j�3����ǟ�u�o�e�d�`�n3ԛ̿b��Y�PG�(C�A<�Z��B�\��G�8�*�# ������a�<^�>�rK�r���a��HlQ/��?HY�S�h���f�w��)�@���*�nӜ��Hǈ)T�u9���3;5��ؙjl.��{
��m	���Ʉ��:�5[�] �4�$F��߽��tQ46- 	Iz~�Gy�'W��	]�	r"Dd���꺖Z(��!�Q���y�,n���w�� ��5�AkTRY]���p��1�����+?��5b��Vu���|/���ϣ[���A�*w!�I��=� I	y5z��<$�W��xl��2g���z`Ε�ھ�i�䰥�R<���Jq���x�t������5���֡�&Y��V��O"�|:�@���*�n���W����]�lEGV`2ɬc��WN<�V�QK�}2r��q
�T�P�y�'�X�6q���D��$B�����o�u�/|�Rc��[�jZ���R\h�(E�4��+5��N��M��q\�!P���b6:Z��c/����1m[�d��%^� r��DI6�<�k�`�?��<�G��-^/�eo�L���hl��h&�.���Fٷ�p"�.��탯;\߰{�P�1|j�:"��8ļ���N}�O̡��Xd!����y�8Tc�A�Gd�o[b*7+���Ã�n�٨"�B���zcF�����ٕ��������R]Y��5��X-M�O��~Ӯ��ȏ��F�[�c�Ĭ	�q9+t�}gm����4M̍���#W2���j�Bd��g\�Ҳ�}�-M�O��~�Ѩ�f?�R��h�	�l:\a�	�+4D@? �z��J*��_?�v��9�2�LX���ֻ�x(�i��/RŻ�&ǥ��a���F�LFC7�5$�)�vx[&ᱲ�������0+C��Q*S� w����o�c�fm�հr��<Н����T(rf�����E���Xyܽ%�J�0�ǻ7t��L��=4���~9�n=*w��>88a�`�f�:3b���qq���"�Ee�6;�c�fm��Ƨe7��
`����0�E>�r�����6?
-9a��&5�/h\Ef�>neb���.�m���=+Nh���/�Ԭ!��Tӧ~\�)�`"���b���g�d��<fϹH%�P�7�f�:3b���qq���"�Ee�6;��\9�oA�K�q��D�7l�"b��"�#�fp�J�!F�R��t���(�x�@�
�����Pع���;Ȼs����~JFNǙ?v���cc�5D��0h\Ef�>�QI�w/ˤ��d9�=>����o<���Hn
V~$\�tj:��sQ頭q�a�[��9�β8�P��G�=4���~9�n=*w��\��N��-M�O��~ӎ;�z��&5�/h\Ef�>�QI�w/ˤ���[6��1�2�w��_3�mE�_s���D+P��LFC7�5$�)�vx����a��2�����Vc2�����Vc2�����Vc�cRq>h�S��P�T��x}W�S.L�t�[Ջ.�ocF���(ZH4~��2�����Vc2�����Vc2�����Vc��G�ZB��'+�3Lَ`�M�(�GO��-b�Zj�����x��Rw54D�����a3��D��Lh������Ց��a��|�� ��u�螔m�l:M�� ��u��?�7
���� f�Lu�m�9�2�L5��_ۑ;��ѥ��,�?�Bd(֮��.���D�+�7�����L~΄gO�3f��*�����R����b