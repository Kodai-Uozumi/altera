��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���a?K���J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-~09h�i�Nq�{5��]�0�lK'���Xw����Q4f����om2�YQ}��1\���^�9:�M��z�}�I@�;摼ڃN\��~�����]��i�i�n/�NE��l�JHn��z��[�Q-�͌4s+�ny����@���_�G��G;5B5Y+�Ȩ�� "�Q��wjw�K؞FMN�*�])������u���B��C�QU��}<o�Y�d�*�K�
���A�F�7���3�GXS����E@��~���($�J.���
�=W�֯�^��N�&��?�2�1p���}������]�0�lK'���Xw��_
�u�m�\��q�Z˻r����4��a�&�������N�N���aC�h�>W����Q�\DR]R�x!���2͖梡���h`�fx*���-the���ʝyzL͊�q��5�?����F�U8�3���lHc�,�u�:��ܣ|4�/��ӝ�9��,V z�J��x�]Ҙp��0c|=}�? ��i�+���9�)bv'.8��>oUa/�OZ�5�p�������m�X��Y�$���e��y~}�;h>xQ)JC�4];ˍH�ƽ��s�I2�}1R$Z�#�u�q8�6K��uIm1��y��/e��^p@f�Ԡn�gg�L�@�1��ꓩ�l;��!I/�������A��1��+�W��J�ݨg4$ _o���6cMH%�]�<o�nïi�;5B5Y+�T�����NF@��u�'�3�$ �#^�Vn�;ۂ��IÙ=�H���0�EѠzM8%�Y~��`�J=�C��a���\�vūx`��:���Ϥk�;��|B}ø��y�w8#�RC�G�G~��6�5�!�7D۸���9��;9k#:̧�	��U;r��Rbˀ�7���E{�ޒ������U��;6(Ӽ�\�v�O$�������:�ʟ�����R�fPذ0������P=mO�u��}�Ӫr�6�����-��w��;�,ZIE)���K�jЌ�N��P9=y���U�q��&�'n�^0o�]�� ��{��j�T��5�M�1�>�w�r�q90��y���8�h��@���Np��['�>+��V���;�z�i�_!gB��L�`���o�C0M���LI���?I)W�F��F�zL͊�q�����x������]�cC��\��z�+�V�&��'Qo�n<�!�A��ؗm��)2��'�al��p=�I�Qf͕vf�'l�2%0��j���c�y�A�
c�M���q��9q{�f��a��{oS�`�]	W�/U�MR��[m���$�(�+
�Ф�kg�ٌ�{m��|�.�=���(��ЙhMJ{/��1!��<U���F��O�uPU��s5�L�R���tŴ���v���~���d�٣��c�A�L'� T囲X���5^��`'&Bc &��L�wR��A�����r�����[�y�95�yG���OI�2+쀡D	�+?�2D�"zL͊�q����)_�����]�cC˸�G�x��7}Ԟ
t�������t���m���
i�kA���8��?��%:T>N,ìp�����o��`z�X��r����Hj�h���89�sfc���r����,n���O����aa�ΐп�hZ63S�݃O�hf>Ŋ Ύ=}j��x=�o�j��\�;��*����	�z�}ݢ{H#�3F�;l�}t���UvI�5U��A����\�v�[��������:�ʟ����Y�"J�p;�j�`,k�M��/��	���G�¨0nE���[I���$M��T�?��w̢��f��׿����8�����p�;ۂ��IÙ=�H�k�0W�)�Q���ʯ�V}..r!��i�>��=h���+ᘱ���#/IHI��F�;9���u�!uqE&.�?��m����z?`�D�.}���N�@|W��W���b�$��Um���s��-���6��z[���"�WT�j
�I��w��,��xc�lL�J*?��	�2�fr1y�r��1�1�WC��nk����Q�Ar+A=?�<O����בa��@IE�U����S8��y�)xʔ�]44�t-��T�\ ��>{O����Z�M*Gg��q�J��G���~����0_���>���̈�1�WC��nk����8/�.���Ҏ��� �E�o����TD��-�`��8�4���H�i���"����3M�b\�-����R���\�TY�[��5��+'}���PI���!�	�������׆��M��li'�8�`�Ii�I���M���d�W���-��w��בa��@IE�U����S8��y�)xʔ�hMJ{/��17�v�ԯ�{Ro�č�tI��6�)`_46C�󈷙�����q��:4\x�\��r�7�v�~������]�!��	Ǹ�y85��3}�@�7	s�A5X�g��U-�eRAѭ������\=�����9H�Y��oy�{�<g�E�.1�u��VD.�+��r�3�C􌇷MV'UK+k�4��r�*%�E�=$�O�夡A�����<��z��}�צ:�)�6�����}כS�]�Jg����-c �ЄW:)�%��2�?�c�č�Y���S�)37J*u�v3���?�N"����y��,2�����^���@�c}-Wh�4�B��ٴ�F6_%v��w\�f@��ͻ�U��J�'1�3��u9j1�f<��z��}�צ:�)�����qZ1~�g]�I���B��&���a�%�j@c�rn7Zմ#&$�ZN�I��+�R���L�H,�jЭ��9�p���e'��ǩ���KT��I_3#ڸZ鎬����b���h�6g��$y�z��eU�e��������Dg��y��tqӴ����s��	�54v��ei�;3��|�QtDo~e۞h�G��L/��!n}y���q���U��Z_�� ���ѡ�e�LZ\^�e���Eы�`�M7Э���j����H��[n��B��X�g^�*����)�%��4_�;��	��L-�yC³��Mz��;��ҋX����0�a1i~J�_�]w��ݏ1��𠛕!��L�ވ���ۭNJ?�s�C�,����e1̙�;`�r��̉'�����.J��h�D��0.�f�;�>)ʡ2F������|��].��'���Xw��Aدo�zea���||��/8'�G~+�3;��\���\��k�zph5)�� �T�5B���"�D<��ͻ�U�ES}�T����3c/��!w=����^<��z��}�צ:�)��������B*�2���u���d���=A�2�S|���f?��� <9�G��7������!�<GO�\��'��o�/��2�K��v�~������]�!�����#e�`�%�]�]�Jg����-c �ЄW:l�mq���)�:�ۇT�0��e�zt�z��Al�q�N����h#!��ҩ5>�����O�D�!n}y���q���U��Q�����p ���ѡ�e�LZ\^�e���Eы�`�M7Э�v�4�oe󕣢�'.F�U�#1Z�'�+k}��eC��曽R/�WQ��9�p���_��cZ2Tv�~������]�!��	Ǹ�y85���~�h�Sü~���U��g��U-�e?�:�Z%Y�uS��ݏ1��𠛕!��L�ޙ�t��O�;>�z�*)=�*c>��3DdZ0o�vʓ��<��Ӭ�t�$�7HfVutְ0�zǵF��^��0� �8k>6s����]�!��	Ǹ�y85���~�h�Sü~���U��g��U-�e?�:�Z%�~kE#z��eU�e��������Ӟj��s �׊�8²u�8���=ON��t*���һfVutְ0����Uw����Ig`i7G#+�Ǵ^:�+�	�t��q{;�]�Jg����-c �ЄW:c��;�&����\��z�+�D��Lh�Q�%Z��;�t.r�����w��������́����H��QU��}<�&���
k:L~΄gO�3f��*����f���,�L��1\���ch& ��I�p\�WB]/�oRA�N��E�EX̭����oP�{���$�r�^K������О.|��	(���N��B�)Y]��Y�,Z�J
_䆼�\�v�<A��s]�(�晅Pt�^ֻ��)�cOKO&8^�=�Q��M:��2��w�怖�č�Y���S�)37J*uc�A�L'�	�Vh�/�owђN�~R�wX�մ7��"�5�č�Y���S�)37J*u)T{6T'��9��tH_3#ڸZ鎬�����G��{�1���=����|��].��'���Xw3vm��&��u9j1�f<��z��}�Q2�+�Y��'\��v�~������]�!��N%��9Cl���&k���!n}y���q���U��=&0�k���Ig`i7G#+�ǟ
��|�6|�+�� VU+I��(�@$.>�~�Ι���H(Ť"Of��3f]Ǎc���L7ܼ^GI��'�,����|#^�Vn�^ֻ����XP����w��$C���2c�'z͌4s+�ny�X��{��ܛ�	��|��	(���zL͊�q����#N��RmHX���2c�'z͌4s+�ny��#_��Y~��`�JKݗZ:���'n�^0o�'�=��d&(C�#�7#^�Vn:�}��E5��*��w
j$8c��� 8�2s�. �͌4s+�ny��d�X7Y'ʯv!	��q{�f��a�:&�>��s��%�a�*k������Q��\���;ۂ��IÙ=�H��^�7^/��=�k2B]p��h$���RA8��'n�^0o���{����I��'�,���<����c���$��;5B5Y+��q	k���A /N��#�D�D@���גy���	>]��|��~�Ӆ"�5͌4s+�ny��d�X7Y�~*��d0�^ֻ����XP��ȁCڮ#�$�|�"Y�(II��'��%ȣ��.�}!��}����H\�iba�G���6(g��9��������HJHn��z���z�O҈LU gZkk��g`�.����?˻D?���W����r�Ch���瀜!���Aq{�f��a�:&�>��s��%�a�e�ٔ�"_��z��"$Y��X�;5B5Y+�T�����N1�*_��h���W����r�Ch���U=h�.�{��)Cs*�t�'n�^0o���{����I��'���Hm~�k����w�,�re��BzL͊�q���`���ˮ�5����`K�0�Dʒ�<�iy�Ǽ��^ֻ����XP���b���DY�9��'E�<lG�"*4��c�����\�vţ��W)�:w͌4s+�ny�|�uwu[7F�r�f�t9�a��j=IÙ=�H�O5�#S-�󕏜9����V)ׅ8�﹈�iq{�f��a�с�'sIP�1�*_��h���W����Cw�Dҡ�y�3�Y�`�'n�^0o��0'�c7�d��Lԗ��|���\j�L�������.G��~Z�7�KXͯ��<�0�Dʒ�<�iy�Ǽ�1�*_��h���r]c��{rϤlΔ^ֻ����XP���N�GU��^ҝ�Ȑ�W=�e+#����?˻D?	���fɻ�n�j�Uo&�Y��>�Z鎬�������(���Ru�A^H	s�A5X�g��U-�ex.u����57�I4 b%�k]�s���D��ޡ�{�50�Vr.W���ۗ^4/��?EMf���9���q���U��F*D@��j��pw��˷���d�φ���;/��.���w��S�[�QTߨ�O3����KCgpzl��a�� �܈~\�Mf���9���q���U�?�����"2�#�>��~���1��B����qC�<��1���?��;���H��Ig`iZ鎬�����7]=k���1�&"i�9�����>l\�}�jT%q�#��]�!���äs_���l�mq��L��T��>�]bU9]M(��۷�_,2Q�U	t�ޯ�l��ljT%q�#��]�!���äs_���l�mq��L��T��>�*%˯S�E��۷�_,2��K�Q(�I�y.͘�=Y��_3L��'9���_�sL�j�赒�^ŇI���FC5��v���ѻ�p�5�e`��9-Y���".7�ﻋ-���L��&��dK>��{�T{0)V�Wx��4�so�	�CR��$>)��8k��t�7P��T��]�!���äs_���l�mq��L��T��>���VuS!ִei�N�iP+�����u�	NMf���9���q���U�?�����"2�#�?�< TL�MT�5B�������;��K�Q�c��Ҏ��=Y��_3L��'9���_�sL�j�赒�^ŇI���O;�2��~��ѻ�p�5�e`��9�*7��x��ﻋ-���L��&��dK>��{�T{0)V�Wx��4��]�R��$>)�0� �<���7P��T��]�!���äs_���l�mq��L��T��>���VuS!ְ����Dj���������	l�l���Ig`iZ鎬������=X�~���X%���xT����"8M���&������Zp y��Pc��?@W�b�$��ŏ{�50�Vr�t�����`�]�)ě����-�$��]�!���1����mӑ!�;�?�R�����Ouܲ�?�t��d�٣�����6>��T����{o����(�G�|F�d�٣�����6>��T����{G;9��Pj������C���=Y��_�@5���<��#Tж��)�f��qb�2kl�
�]�$��'���Xwa'�<� \�_Q路��+�W��h[���� ��ﻋ-��� 
���u���ۖ�lh�_�s����^E��fi���K�Q�R��9�u�!J�ǂ'��=Y��_�0z�cUL�ȘB�k�^ǙPn�O����	a(􆿳���t�$��йt�����w�$J���Mf���9��Y�{'%sgeߪ�{�x�#!b�PǨ�o*� 7�v�ԯ�o��f�kѶ���� N�B.D��z��a7��ﻋ-��� 
���ua�4f�+��ۇ�o]|M���k Uz�Q|M��K�Q�5����`K�WF��0g���~��n�'���Xw�j�7������i��9�#����c�T�\ ��R��r��)}���/�	q@��57�1ʾ�!�������Y�Y�{'%sgeߪ�{ޒ������JoEѰ�MM
��,=�*���BQU'�����p�m~|��^�����K�Q�5����`K�/���������D����'���Xw�j�7������i��9�#����c�T�\ ��퍥6�u!�y�2ۆiq�L����o�>�5�ﻋ-��� 
���u�z)z;%Ψ�w�Ua���+C��5|M���k��s�KT�����bpj��6ג�������XSx�lޞ��rs�i��ߖ� ����[Ѱ�^d7�v�ԯ�o��f������bpśL���>AU!"k�Sx�lޞ��rs�i��ߖ� ���y�:�B�)u�%N�ߌNu�5=��a'�<� \�j����fX)��F��Y�W�x�D�:`��nZ鎬�������(����YZ��,��<�^0�h���oMM
��,=�|.�Tӏ��U�^���OV��6�� ����˭b� �X�Ԩ�d�٣�����6>��~u!�3Vt���so��㸒�ﻋ-���C�M��N�۔�Zr�X�ȀY;+�z�;0��r�0X�Z鎬����Y�V��#q��U�^���ך;�gP�m3��>*����^�'���Xwa'�<� \�j����f{Ұ�f�>��֑xGV��hΤ�`�ό���.���K�Q�&������(N\�(e\`�?g������ݘq���U�pzl��a��m�6zi�(�O�%6�m�±��m|���.
Tg�ﻋ-���C�M��N�۔�Zr���)�b�To��(�D��=Y��_Q2�+�Y������bp�N�|�!������<��!����]�!���1����m�6/z��q�lN}Ot�z��a7���d�٣���$�j���&�Y5U�R\� �n::LF�a�{�50�Vr�؊�"�D�3l���|g����A�e�]�!���1����m���Z3��Z{1@.&��kD�C��Z鎬�������(���x����T�)u�%N�ߌNu�5=��a'�<� \�nP����H0;��eݰdo�Y�ﻋ-�����S8��/C��kX�{[���G��>ٮ����l%鯅��? oOB�Cje����H$�DZ� C�C�.�.�;F�v�f1۴��j�n�qW&�]�ר�]�!�������͋���g_��mQ3��T�L�L�`���������"sYwvQ-��̡��Xd!����y�8T28]��:�q�����NF*��_?�v��B�>�9�d�٣���9�����6�<���sW��	]�	2�n��tR��s��d�\��MN����!I/�������A��X�@�5��6�l��sХ+�:R 8*�A��jeN�V�����׷eh��S��L�u�RmHX����20)�_!�D̯k"a)�m�d�so�}a�C�ub;�;��$��ľ$�o��>
��a��Ls��喐Hj�Y�_�]	5�e� $p\�>���S�w҄�|5��s�#��v@���J֭��|�����]�Kt�E*�#�,���ns)��E�$�v����ox3��vC��Z�G�a}Cy^6gVW���%@�~��e�0����5Je�4o�}a�C�J;����t�A!�?7L�sZ�	Tt$�ْ�6�j7 ��Lc�TH������7��ZΪm�T˚�Jz�0���je�Vmf��}S���u�����!�.3հjdo59
4/�]��	�`М��Wa;@��{�;F�~��j�q9t2�����Vc2�����Vcl��w&� ��tF��J�[��<X�����Fu)n2�����Vc2�����Vc<T�R�$�P���������$OkY�Wm���Ժ	<B��g�9y�>n����"W���P!��|���ř[�~ݶU���[W~L��?�Tm#����Xb�r�I �۞h�G���',�K/{J }dx>3-���t�q9캧xӍ.�����{�T�ؼ�n�B�'��D�Mp�=n�٠��f�;�>)��-oO$t�&k��@f�6��	=Q+�����3c/��!�����g*�s��I�-����캧xӍ.�F�Y�H�n�,�E{�n���
�`}����`w]�u��;�H���o�Iy��A�-��N����u8ۯ�p�O��{��f�;�>)�,Զ�1�J-��N����u8ۯ	����۞h�G�#�2�����,��f��=H���A��2�����Vc2�����Vc2�����Vc�ǑW�A Pc��?@W�ȎY�I������[�,�B2�����Vc2�����Vc2�����Vc~�<>�TE`�]�)ě��;��K�"��-�y�T��\O)%���J��5�P3 C��;��K�"��-�y�b��:��e|��]to��񐙣#��U	8	EZ2]�oڭT��ե�o� ���ݔ�H;"�g~����X,�;ڒ�!_m���_A9N��b��ؚ���$��k���I�`?���d�2�كs_����fB_D��h>���ih%���J�Z(�1O<�I��.�{�)Ʒ.���D��u�w�D�{xH:������Æ��2�����Vc2�����Vc2�����Vc2�����Vc�m7���ew�՘��nIDn'��Ci�Ed-� �HB���$V2�����Vc2�����Vc2�����Vc2�����Vcu�SgJ��V��Y��/���o�v�Gf��(�;����{`�*���Q`P��^���\�}�����	���9W�z~�Gy�'����KCg^�n��UhҢ���I����BUt�a�ke[��u��}�l�1�����0���!�T�.�O�[�]���4�磕���ɞ��C�g�0�u��a�֧�I��3��a���	)Ԭ�>@X��WG ��Z$R�Z�]�+u�CX�N�g�c�`�N�����Å���E���#H��b:�N�NL��,��u���R��	0ڳķ�;��|a�&3f��t��U��$�K���6f� 9{�P�1|]6�>����U��\JDR\�=φܓX�H�->t��w#o�]�ʄ�"�G~4���t���(�x�H��	W��N�g�c�`�N�����Å���Eۃ=�0J���x(�[.o�;n3�#���۵\��rw�&�z<aSm�6��`4�04�jf��ܐ�}��JdT1�V��	��y ���l���L��k'
����1�a����KӴ��^�=� �9D^�����i�ê1iKS,
_��s�֙f����hڜ=E��r���qb�H��j�s�jd���lj�Ï��	j�ە�((Ut�\����'|b<���1��X��WG ��ʙ���2e���T��?o[v<�F>��a���!��G_	���`Xg?�вp�cA�	s�A5X�g��U-�e��$sb���x����u���oVl�(�!�G}��z��9;�B�|���qbsZ��"�)�{�°!�?����S�)V��B�1%�x �N�t&����1〈)�����d��-��!rϚ����5�P3 C��Pع���a�	�+4D@���'9tT4]d���z�'r�_�(p��ӎ��������Ս*�(f�Kp�-a�D͢fU�9�׏�����MFi��|��wØ�ߜ���,�ǰH7"LTftpϣ�و���G>a%�r�����>��Z?�7�!`��&Y��V��� �1
e�UѦ��	}p�m~|��Q�7��UO/D�;E���h�}l���L�C���ea�Xi��Ԛ��b�$*�&�P�2�P�L��M����z��R�rb�񄐙�#o�]�ʄ�"�G~4��X+-U�9sz��c� �-M�O��~�n
s�] ��z�S�Lw΄�WV�����x(�[.��T��?Bo��ޯ��k=2.�4��Ɲ&�K���L���4�04�jfx(�i��/R�*�W�Ǹ!2�͞nOY�����	���9W�<�V�QK�}����{G;]�jz�X�}_�nx��?�uUn����:���|cKE#�i閸*�FS����Àgڿ[�F�}	��x<�&Y��V���g����/�4\y��<�vd�̪�Vx����NӶ4[k��#D?��HԮg�~3���ix	�"�"�5����`K�Ia����y$!Z�ni�A|'��ci�]�N	�!����l�z6r?�1��	�gc��`c�����U+t�+����(v�����1nE����y=�~�(� ��*"����[�����#�A���k3���s��Ö�^��iHP�k~��>hE���q�*'���%G�	r�w���W��.���!F�5��!��G_	��4���_�bR�QP5�E���E���V'/Ρ����qt� ��p��F|�����_������%��[� �����CO|2�@xZ@4�׻��Ƭd�e�Y���T�+Z;1�!S)%ۆiq�LԵ�_չ�ŉ��7Tj)��0Y d��`�1v�-�/D�|11�Ĵ��j�n�q�9�2�L�5����`K������D��C���,��Lq�"��2�Gq��	��0a���ta�a�~vT���_���\{��x�gL F��j��H0;��e�5��[K�@���'R���#}ؐS����Uh1�b_X�XV�b�z'hۉ)��R���+���Ã'�� ��,�`�]�)ě���7�����g�0�u�7�b��`�]�)ě��Pع�����)�l�l��E��႓ߛK���8�z��c� �-M�O��~�e�7�L����w�a��D ML:�}q^J=����\n0�8�;������@ګKƂQ��x:A4b��JB䶓������Ut�\�j��ӏ��t	�,^)�%�]��8��w���>-�F`z�k��h m<���HK���b�([��}qn
V~$e�7�L����w�a��D ML:�/�}q���V�y�Gr��w�a��D ML:ޅ��J���J�1���K���L���4�04�jfx(�i��/R�*�W�Ǹc���2�@ �"���ʫ�>��E�>�oR"�pR���	���FyL�&��8]�]p扦�2�0��a(Qݞl;U��+� ��_ߺ��5g�)|���:χ���^ǙPnw	"�d�kL�|Z� ��_ߺ��5g�)|���:χ���^ǙPn`B]z(,� �ҋ�;�0cp�h9�c��� � �9D^�W����,��h.3I�;��|B���%���lq&�3�N�0��B$r�Ch���U=h�.�{X����O��	�����Q��m�J�
�M�٥P5���rs�i�Ǘ$� ��������,%�ۧ�A�YQ�(�O��Q�����gV��|���\j�<lG�"*x�©���P*ra*�٥P5���rs�i��s�٭�������p^�i1_���I7��-5!L(��̭�`����2lq&�3��?D���Ø��t�Y�x�(!M����A���gq�$dШQ;�im��|�L�݋r\sQQF�;�?2^�9<o�nïi��ٛ ?+d&(C�#�7#^�Vn>�1�1��_�G��Gc��ҭ��^ǙPn�)�����\���9�}\#�`ށ���y�{�'$�7g�@$>�	}o2�1.�@�Ȼ-�v���B$~E��sp֟kh��=�er߮�fӥF��򴖇��/��~q�e��ͱ_��Yu��Ǌ"�x���|���3U(�{Hl��O����	a(􆿳����	S��7��"�5h���X �Z�^6ː��h���X ��f�;�>)�i���F�}?��qW��nf|FN�7�gI����I�}jf��k�-sjv�����P��
���A�0sFw�K@4I_�GZ6�L�25�%l��7O�3 ��f�;�>)��gH}G'W��j=/x9�=�Da���B������@.�>�ȼWt�MoSN���ˎ.�1������yA�B"�u�������D��H��u0޶��>_$;��|B4Y-<L'��s��;��NcQx�Ԏi���QQ�W��vw<&?������Z���Q��m�Ү����,j�W�q�l0���2�W�ub���<p�ve�}��i�Ɣi�����Q�@�p�~ge?�΄x�g��	��S8�t޶�2�z�`�0+�O����	扦�2�0<�iy�Ǽ��Y���҇ct�:��RE��|���\joU��՗7rx�©���P*ra*�٥P5���rs�i��T�ۿ�#�dWp(�, �dh��X+)%`d�Y�8!�iIp�2r�o�#7�cL���	Ǹ�y85��3}�@�7R�����3U(�{Hl�3��rm��<�䛄�� �f��K�S�U5�f4����;>�P=��J�xsEqFM�ϸ���K�ْl��]�B/��v
���3ľ�Yx�<@���U@���:��F��L{����t���6��^hq��:�����]��Y�,0��������a�̏���eh1q�c���	?���ֽ݅u�x���|����G��8n�$�؁��ryO#��!�!]���px�y�;����&��0�m�4%=3���!7y�x�~h�E�  ͎��7�o�_���p�*_�uFsY�w碆�����<`��S�v��eh1q�c���	?���ֽ݅u�x���|����G��8n��O����	a(􆿳����	S��7��"�5h���X �Z�^6ː��h���X ��f�;�>)�i���F�}?��qW��nf|FN�7�gI����I�}jf��k�-sjv�����P��
���A�0sFw�K@4I_�GZ6�L�25�%l��7O�3 ��f�;�>)��gH}G'W��j=/x9�=�Da���B������@.�>�ȼWt�MoSN���ˎ.�1������yA�B"�u�������D��H��u0޶��>_$;��|B.Y�X�"��6j�"Hs��S�<뒯2�����Vc2�����Vc��Y7�N����h�^'��_<V[HB���$V2�����Vc2�����Vc�cRq>hM?�(�v��s����쪄9C���8������V�2+쀡D	���me*;��|Ba��M(��霱�"��7����)�YCHdpQ�8��+�:�ik��+ņ\.~Jc��z0��mWD��������G�C׋	�Kv�ƞ�qx�����tÎ$*V�����-��A��D�V|�)e����ǉ"h�%��R���>e#M��T�t�mQ3��T��{<"�]I��=� F��v_}`_���~�̒���Ue�s�z�:�y�g��}A,K�-��_�U qKj;M꩏�D��#�u�q8�p�m�If����T~����1�fT_UXe�̔��?eM�k	�xw�<2%�	�}:{u� Q������L�C���ea�Xi��o����Ӫ� Q�����([��}qn
V~$�d�?�4��2��� ��1��J�b�z'hۉ)��R���T۳�͕���?�I���6\�4�@���(�?<-M�O��~��D�$0�<����5>!\��쾋H;"�g~����Xz��c� �-M�O��~�/tyc�����>�z���	x=:���r���9��j��6ג�n؞�
�WW<����,0=]^	�&����ג��X�H��C�j�7jv�]���r"nCo=7�}|��	��a-6�Da�d�?�4��2��� L޹��Q&��>�z����/����٥P5���rs�i�� ;O}�I:�K�Rz�X
3kZ��5ߧE4��n��kc����d��,�XXuUt^�{�Kو��. W��pG���9��,�-�0�,U2@x����O\��؂��y'��BS
��T�Ch�oCL&�x�GR�ø��-�jr�*k�������:���d�h⎙l�� �:w���9L��ѧ�#r�#AXӾ�T6e<�vVҹ���Bo���+���|Ai@,��yګ?�����DX��`aU7J��,��{��X j�*�~n�$�����Ę��(8� �G���0�����F'�Z��%g�|m�$a�������V�¹W�`� �h7 �J#��X j�*�Mx<�IJŤE���!�9�Grw�&�z<aSm�6��`4�04�jf��ܐ�}ļ�®���Aj�X���{}�=�v����KCgDV,�ـ��+�`4�M �m�`h",K�-��_��2$6�sI�f^��h%O��f]�f��%�'���B��ôZ�v�~��	�� <����X6b^�Rt��Z�)�Z�(&)~U��r��3K�[�·��`4�bi����͞N	���IyX��,����W���l���L��k/���`D����	�W��ٕ����ޒ������y�N� Kp;��|B�M%>Y%�Μ=E��r����%��֊�0h�5e���a�֧�I��3��a���	)Ԭ�>@X��WG ��Ѩ�f?�R�����bP��a�	�Z���o��񐙣#�S�T��=7�}|��	��a-6�Da�d�?�4��Ӵ�"�6j��7��|�K�U#:�SD���s ��,�Y��?�/����s@L�Zao�o����Q�?t�R_�f�Hى��_�
k\�^�sW�w��fD���򫒡�W<�׏�����Mrw�&�z<aSm�6��`߸��S�Ȍ�>>Y�k9;��|Br:�j�@�s3����َh�D����ŕ��9�z��o2m�-�Ce-X��y�:�B�{�@�y��?�d���&��d��L_�xw�<2%�a�ЗU���HU�:=�m�`'��<��Ȝx�� BN1l�n
V~$�i��"u��H;"�g~����Xz��c� ���,�^'t���@��T��R��a�J��vT����}�o@��ѽ��J�����V%_�E:b��Ut�\�m�O�����(����jq.�w'-���J8BW�R7�2ȰTl��W ���t�F�fy�o���8���~կ�}�aá���(�^�G���=�ni[�b��o�CHn
V~$(|��s�i�OV��6��:�j����y�ٛs��1^~�8���d�������p^�V]��}-��\4v�@���rahF��v_}�bE��`W��U�n��*�%�UL�Zɒq�$�P�D��P�����
��M+;��|B�&byG�O�˵��[�x(�i��/R#k�˟ܒ�o|k�Lb��ܐ�}��JdT1�V��	��y ���Aj�X��룄���~�b�Ƹa���IC���U�"�510�p)'�8ϳ�po��z��X�j�{~ �:}#���3a�.��Ǌ��i�ъ������&�!+5�13"���e������.�G�����so�:�L���l����/Z`�k1��r��Mڼ��:Q�@z�PS�����b��T�Q5�ŁG&y�A&�/)��� t��]�kj�U�f��&������̑�z���t�P�'�6�9���gbc��� �/?z2�����͋�V��Ĵj�O�&�v�3*�ԟZ�S�h����� ����΋�
,`mu��.8�&�������^���<�o�2JC�j%�~R�`Z���>.?��.7��Ŵ#����#g�k��m�O���rd�d�JR'b�'=�(����`Q�f����*d�����}�o@��ѽ��J|�����!m�O����dQz^Oыq�GR�/!�f�u�R�����O-���8ǻ�d�?�4���(�O�%6�m�±��m|Z���Q�K�]��7�0�/��~�j<�ڦ�`��B��������oP9����,�ǰH7"LTftYD3���L�%`�/���@�Wu�t�Ru�A^HG9�Xb�P:�WV�#a؄�Ș�-U���4�磕G��64�kG;9��Pjs��r�F�Q�bc�+�(��?c�O�F�Tr�f��4i�׿��/v�R*E���&�Ut�\��d�?�4��Ǌ��i�ъ����%��v��/tyc����(t-�D��ht��g��倉r˲����x�ԉ�>�&�(5�;2��dc�@z�ׅ�ؘ��N�g�c�`�9�d�L�B����.� \6��.Ƨ���bP��!���2�(/ѿ�����Q�9_*p4�-�C��7u#md��X+-U�9sI�ߋ�N�g�c�`��L�ΪA���-�廈���R������@��bS���+��-M�O��~��6��X�X�ȀY;+�z�;0��`����n'٥��gV�?5'[�鳒��@��T��R��a���3,ő��Hp9��T۳�͕��/tyc�������so��C$WE���z��*�m���ɛ�?ө(|��s�i���R������@��b�x�. ��#P�j2E�?�5ߧE4��>je`��@d:�����{~�&�������y`Z�b;��t�o�� �-u���kn��8>��LP�,{ω��5`����!**�w���!X�uA���|�wƄ�{Ƨ\L���jߓ�U��Y���zU�J�������A�H�f-�M��������d�?�4��[;T�!'ؔsy1�n��뾦�c�}���Fo|k�Lbx(�i��/RŻ�&ǥ��4�����-%��ʦ0m�O���{Ұ�f�>��֑xGV��Ee6���uo�Mj:F�S��/�j�LY'�P�h<���8-I����c���1�ā���"�1�C���N-�y�;�a�ke[��u��}�l�1�����0������Yxkx U�_@+���Ã'�� ��,�C�����෨J	a�ЗU���HU�:=�m����y�BDG;9��Pjs��r�F([��}qn
V~$m�O���rd�d�JR'b�'=�(�q9+t�}=��Ez�wq=0�>\�(?i˸3�J�
�M�'٥��gV�m�O������W2���ݟ=�NM���ɛ�?ө�&�(5�;2��dc�@z�ׅ�ؘ��N�g�c�`�9�d�L�B����.� \6��.Ƨ���bP��!���2�(/ѿ�����Q�9_*p4�-�C��7u#md��X+-U�9sI�ߋ�N�g�c�`��L�ΪA���-�廈���R������@��bS���+��-M�O��~��6��X�q=0�>\�(?i˸3�J�
�MɂMv!���x��a�z6���-�廈��j����FA�$����@/��r ��%�z�J���d�?�4��[;T�!'ؔsy1�n��뾦�3t���=�4�04�jf?5'[��jv�]��a����g��a����q=0�>\�(?i˸3���I����?5'[����s\������N=�m�6ziǊ��i�~	��}q8BW�R7���r_��m�d�?�4���W���2ȼ�mˊ��դ�Hp9���d�?�4��Ǌ��i�ъ�����e���\���rK�&���&S��"��hTC�G�L奟gke�(ƚ�4j�}�������A��(/4��]G@��z"B�4��X�q�hH0��^o��[�u`���ҕ<(�(m�O����dQz^Oыq�GR�'�^�����P�HS|�4�04�jfJ�1����ݾ-/�φ��<�6�)�@����(|��s�i�nRdd�����C1zh�I�V.��S^~ߝ��wh���t��d��WԶ%T��Cz�A�uG���G�Ȧj��v������^�n��Uh'��x�-ڄzI������j%�~R�`Z���>.?��.7��T�$����Z���삕�Յ�.rV֡�{���F���B
lE����7���� N��r*Ѩ�f?�R�^�*�ǒړ��Q .�L��H��	W��N�g�c�`/tyc����s��1^~Ϩ<Z.َ�>�1O�ME�g�������(ӈ��Z��&61�e��@F�KD�Vr[?z%CS2b�ү�+ҋ�K:+>��-�廈�OV��6�� ����˭b� �X�Ԩ��1��X��WG ��?5'[�鳥����N��qs�@�tͱ_[��nF���<�W�.�P��c3რe��@<����5>0��d����v���-x�@y��.'��w������"�2�C�� YI�ߋ�N�g�c�`�6��X�W����<MN2��΢g	nܵ,��L޹��Q&��s��1^~Ϩ<Z.َ�>�1O�MN�*���~_Z鎬�������(����૙v�2�>d�ܡ�0�$.N��p�-a�D͢G^��w�x(�i��/RŻ�&ǥ��4����K}ͅh�K]�9k�
"�śL��ł��p|3�ޝv�@��s�T��P���g�0�u�?�I���śL��ł��p|3�ޝv�@��s�����Ja�vݝh�c�A�L'���搪zW������p���?���`�te� �Ћ�3���ү�+ҋ=��Ez�wX�ȀY;+�z�;0��`����n'٥��gV�T۳�͕��(|��s�i�nRdd�������O�g&xdp��K���L���4�04�jf&ظ�����C�j�7�����N��qs�@�tͱ_[�+�9-�i"'���Xw�j�7����}�l�1 ?�Ia�f����Sl�2�>d�ܡ���u��X��WG ��(|��s�i���R������@��b�x�. ��N�SF�eśL��ł��p|3�ޝv�@��s'���'٥��gV�T۳�͕��(|��s�i���R������@��b_їE���N�SF�eśL��ł��p|3�ޝv�@��s'��싂Mv!���xx(�i��/RŻ�&ǥ��4�����eVH��HX�ȀY;2deM�|�'\��i���w �w�d�?�4���T^����4D���tN	L4u����]�����;��|B��}H	��*Aj�X��낭[n�_��b��T�Q5�����-VL�ސ������A��(��o0��X��@�v�ٛ�S�a�nRdd���`����n���1v�C�� Y�i���>oX�ȀY;+�z�;0��E'	���M��1WzX+-U�9s�i���>oX�ȀY;2deM�|�V�H�N,������	��c�k�A�(�@3l|�gV��r+e���ٿL��'�6��^,�$�{'���d�MjW�Ne��F�2�C�T\j�� ��������{�H@@y�t`��tH�v���-x�@y��.'�!�w[�/��~�j<�ڦ�`����;dנ���D-'��7gz^N�W����Rg����%�����	�ʉ!�S9{Ȝ��@�^�n��UhҢ���I\Ef�>���b"�r��4�9 I�������p�<�2�Ҧ1���Z��(|��s�iqh�e��+��9�2�L�4�	��m��.��B�����,�ǰN����;^�n��UhY�����Ca�zI�����������D�
���
?�-�Ce-X��y�:�B��K0ю�h;��|B@͐Ov�bq�lN}Ot�l�1C��(��m�6ziӴ�"�6j��y��m�0����,�ǰN����;��e���W�\Ef�>�6����`�}�2���w�xo�Am��uJ"\T}2����؇�8������-VL#s?J�?�{��B�.�kB�a}GFD|`�ht��3i�Y
�,�m�6zi2��� t�&���'H0;��e��Q$ N� �9D^�I:�K�R�q��G��M*����9�!�T�.�xkx U�_@+���Ã'�� ��,�`�]�)ě�<P�]zEW�E��႓ߛK���8�p/H]K�_%�0h�5e��7�b��`�]�)ě��Pع�����)�l�l��E��႓ߛK���8�z��c� �-M�O��~�T�+rJ}?I|`�ht��32O!j����xE<B��)u�%N����Cҷ��e��nF���<�W�.�P��c3��6/�%��Ѩ�f?�R����_��
�Q�Xn�)��d��X��WG ���D�$0�{���F���B
lE���Pع���a�	�+4D@h�Qf�#t�,��r��WdM4@ȂP�U�P���$��"a(􆿳�p;E#M|v|`�ht��3�'�*����$��"a(􆿳�e�&���6rw�&�z<a��r����5ߧE4��p�-a�D͢fU�9�$�)�vxhXY�0
�J�k�n����k]m����
wc�{[���G��>ٮ����l�jV���C����*1^�rs�(�̴Y�{'%sgeߪ�{s��i�y��M*����9���%5�MV�,e�׀4޹�G�Ȧj��v�������k:�(�.��촔��_��:����ٕ����WW<����YU�oY^�h�M*����9�!�T�.�xkx U�_@+���Ã'�� ��,�`�]�)ě�<P�]zEW�E��႓ߛK���8�p/H]K�_%�0h�5e��7�b��`�]�)ě��Pع�����)�l�l��E��႓ߛK���8�z��c� �-M�O��~�T�+rJ}?I|`�ht��32O!j��Љ�1��J�b�z'hۉ)��R��삚 �{��{�9�d�L����{���I�q����.Z�2{4x{^4��*m��L�ΪA����w~���Q��ٹ[I�IT���Va�ir��=Ȣ��~@/��r ��%�z�J���U��ǣB�Z{1@.&�~�����
��`)����k]m��h��7?���?eY��5�g��U-�eԺ=���]�J�1��씑�:��KY׏�����Mrw�&�z<aSm�6��`߸��S�Ȍ�>>Y�k9;��|Bb�lҏ�e6����lG�_�.p����P�f ��ME)��ƽ��Ү����,j�W�q�l����K��֍�`n�P�f;[���w��1������U	U�O� �9D^��쫧ʦ~.���"*��WV�#aؑm��Q�{8���5g�)|���:χ���^ǙPnw	"�d�kL�|Z�%J�bb��|V��	��y��c@�13�F0���	�c`��g�D����E�#?�`�/�vw<&?������Z���Q��m�Ү����,j�W�q�l���M�a�+?�r��Q'�^����m1�H��ۗp���xV���Q����Rz&!Y�Xj՛�֚g���<�H���[��c�Z�~�KO>���͙� �߈ٕ����8�ũH������{�?�d���&�M�߾ol����Rz&!Y�Xj՛���z��"��
��� �����D�2h���2Z�/؈ъp��6?����H��efm�0z�cUL���ޤ�Y5�x�#!b�PǨ�o*� 5���Bi���eh1q�c���	?���ֽ݅u�x���|���N�;5�W��!#���.�h��&r��rs�(�̴Y�{'%sAX���	q�!��ӋD�<qJ�A	D�0��E|�,�8!�iIp�2r�o�#7�cL���	Ǹ�y85��3}�@�7R�����3U(�{Hl�3��rm��<�䛄�� �f��K�S�U5�f4����;>�P=��J�xsEqFM�ϸ���K�ْl��]�B/��v
���3ľ�Yx�<@���U@���:��F��L{����t���6��^hq��:�����]��Y�,0��������a�̏���eh1q�c���	?���ֽ݅u�x���|���N�;5�W$�؁��ryO#��!�!]���px�y�;����&��0�m�4%=3���!7y�x�~h�E�  ͎��7�o�_���p�*_�uFsY�w碆�����<`��S�v��eh1q�c���	?���ֽ݅u�x���|���N�;5�W�O����	a(􆿳����	S��7��"�5h���X �Z�^6ː��h���X ��f�;�>)�i���F�}?��qW��nf|FN�7�gI����I�}jf��k�-sjv�����P��
���A�0sFw�K@4I_�GZ6�L�25�%l��7O�3 ��f�;�>)��gH}G'W��j=/x9�=�Da���B������@.�>�ȼWt�MoSN���ˎ.�1������yA�B"�u�������D��H��u0�۪	�}a?�d���&��w�Pt.�R�j%�~R�`,TK�=_��'_|���;��Qz�#g�k���FyL�&��8]�]p扦�2�0O��m۩���
�����1f���C}���7��6זW���O�[a�vݝh�c�A�L'i��R>��$z����G��8n�3��rm��<�䛄���rs�(�̴Y�{'%sAX���	q�!��ӋD�<qJ�A	D�0��E|�,�8!�iIp�2r�o�#7�cL���	Ǹ�y85��3}�@�7R�����3U(�{Hl�3��rm��<�䛄�� �f��K�S�U5�f4����;>�P=��J�xsEqFM�ϸ���K�ْl��]�B/��v
���3ľ�Yx�<@���U@���:��F��L{����t���6��^hq��:�����]��Y�,0��������a�̏���eh1q�c���	?���ֽ݅u�x���|���N�;5�W�)����P��҇����b���`ܰ��y�{�'$�7g�@$>�	}o2�1.�@�Ȼ-�v���B$~E��sp֟kh��=�er߮�fӥF��򴖇��/��~q�e��ͱ_��Yu��Ǌ"�x���|���3U(�{Hl��)����V!�"M�t�$X4P��Đ/�*�<�>#����*��T����Nu�5=�ò�ˎ.�1�f�8>fd��#���h������b\��7�gI��h"r��f��k�-���D�Lh���X ��f�;�>)�!�#䶜������S�*(�L�U�m�T��Qk��<�o�F�����h4c�H��Y�5}٨5�X��o=��i�h"r����SX�c�,�[`�Oʕ3>x�?8k�{��h�!��ZB4���j���5XsGfh���X �t9��\��9)S.����D�nR�����,�ǰ�����N�C�c���1�ā���N�1�� ��2�����Vc2�����Vc2�����VcREBR�hHr����� ���)Ry���(�䏓O(�e�C�$2�����Vc2�����Vc2�����Vc2�����VcH/5G}}H�T ������Jq��Q�[�AI�Y;�/�4�af�>�4�Fr�Ճ��[�&2����ȥ!Rc&FgŁT��
~�O*��z������n�����ݴV%�Ȣŏ?��!�&�k:����R".�����''µ���XIs���K�P8ٳ���� �d��6=�#�����?t{�P�1|�aԓT�4�t��`�ݓ6+��c}Ex�#Tp3�[1���`�D��M�`;$�l���
F�P?]��0֮�.��Z�H%�nXZh��\���g�nƣ{��!�wd??C�a�)�بf)ӌ���:�Ym����Q~�LL���8�[OJ�k��I�lC����������@�f=H���w/4v6N�'�|��e�q�9	���Usj1n���
V�W�z~�Gy�'��Aɘ%T�T+ ������''µ��y���_Jz������D��ܒ�����[4�����{�`��z ��pOz�$�酻�����塺&Y��V�ɬc��WN :��W>}�s/�]��/��D=,Ϩ4�@a
�l[�hU���r�4�B��ٴ����q6q�^%��=xF	����|�H��6Xw2��j$�@���,-�%�-�/|�w����0�(#;���[|��w����?6z�Y�PG�(�t���C�F�5d���ɱ=��CJ�UF�����dR��:�b��uZ2u���4�磕�}�_�#�ޓ��-�!��Tӧ~������}$@/��r �9���,���n�/������40N�J��7R_'�hs�&o�� 5(Q�g�+%�&;�Gg�d���z��R���F"=�0R*E���&�Ut�\�q쳚�=��v��V�pb�ڙ��Hp�-a�D͢fU�9�׏�����Mx(�i��/R�������a�U�ے
pϣ�و��'sؓ���|᧐���+�|H镊��Q��D��o�Pc��?@W�Օ��t{rо��`�]�)ě�<P�]zEW��ѽ��J��D珞K����dB�4��r����t9��\��5G?�gJi��e���W�\Ef�>neb���.�m���=+��A\/i��KX��iko����Ӫ� Q�����([��}qn
V~$�x2�:��N�B.D��o}����ĳ�e��@���"�2�C�� Yz��c� ��*��؁�T^����H��	W��N�g�c�`�4�!���5(�\����΁�4����_eD�_�*�`3�Z��R P�*��_?�v��[��9���5ߧE4��Fi��|��wØ����Q>�^2�����Vc2�����Vc�cRq>hh����d���]���<в}���hr���2�����Vc2�����Vc2�����Vc��G�ZB�d���nы{��O���u�5=.@%���>ߔth���Pc��?@W��֥��԰{k�2�~���*=p�:���k�K�*��M���5^s�ǫ�����@�ą�.rV֡��@.���g�0�u��y�k���1��X��WG ��Vܠn.� ���6���c�Z�~�ȴ��A�v�i�a����w��ΊB>���<���Hn
V~$�7�b��`�]�)ě��Pع���a�	�+4D@�r�LH'�`�3l���|gݟ=�NM���x�ԉ�>�&�(5�;2
�M�j�����[s������s�Mq@/��r �a�<d���T�����݄����Mv!���xx(�i��/RŻ�&ǥ��a���F�LFC7�5$�)�vxˡO��]�{b�����iLPm�/���?ܸ��Vì�����$(M��AH���BT�^��a(􆿳�F#!�i��J�k�n����k]m�����O��_2��VU(��z�j�L&fL0