library verilog;
use verilog.vl_types.all;
entity stratixiigx_hssi_transmitter is
    generic(
        allow_polarity_inversion: string  := "false";
        channel_bonding : string  := "none";
        channel_number  : integer := 0;
        channel_width   : integer := 8;
        disable_ph_low_latency_mode: string  := "false";
        disparity_mode  : string  := "none";
        divider_refclk_select_pll_fast_clk0: string  := "true";
        dprio_mode      : string  := "none";
        elec_idle_delay : integer := 5;
        enable_bit_reversal: string  := "false";
        enable_idle_selection: string  := "false";
        enable_symbol_swap: string  := "false";
        enable_reverse_parallel_loopback: string  := "false";
        enable_reverse_serial_loopback: string  := "false";
        enable_self_test_mode: string  := "false";
        enc_8b_10b_compatibility_mode: string  := "true";
        enc_8b_10b_mode : string  := "none";
        force_echar     : string  := "false";
        force_kchar     : string  := "false";
        low_speed_test_select: integer := 0;
        prbs_all_one_detect: string  := "false";
        protocol_hint   : string  := "basic";
        refclk_divide_by: integer := 1;
        refclk_select   : string  := "local";
        reset_clock_output_during_digital_reset: string  := "false";
        rxdetect_ctrl   : integer := 0;
        self_test_mode  : string  := "incremental";
        serializer_clk_select: string  := "local";
        transmit_protocol: string  := "basic";
        use_double_data_mode: string  := "false";
        use_serializer_double_data_mode: string  := "false";
        wr_clk_mux_select: string  := "CORE_CLK";
        vod_selection   : integer := 0;
        enable_slew_rate: string  := "false";
        preemp_tap_1    : integer := 0;
        preemp_tap_2    : integer := 0;
        preemp_pretap   : integer := 0;
        preemp_tap_2_inv: string  := "false";
        preemp_pretap_inv: string  := "false";
        termination     : string  := "OCT_100_OHMS";
        dprio_config_mode: integer := 0;
        dprio_width     : integer := 100;
        use_termvoltage_signal: string  := "true";
        common_mode     : string  := "0.6V";
        analog_power    : string  := "1.5V";
        allow_vco_bypass: string  := "false";
        enable_phfifo_bypass: string  := "false";
        \DPRIO_CHANNEL_INTERFACE_BIT\: integer := 4;
        tcd_para_clk_divide_by_2_select: string  := "false"
    );
    port(
        analogreset     : in     vl_logic;
        analogx4fastrefclk: in     vl_logic;
        analogx4refclk  : in     vl_logic;
        analogx8fastrefclk: in     vl_logic;
        analogx8refclk  : in     vl_logic;
        coreclk         : in     vl_logic;
        ctrlenable      : in     vl_logic_vector;
        datain          : in     vl_logic_vector;
        datainfull      : in     vl_logic_vector(43 downto 0);
        detectrxloop    : in     vl_logic;
        detectrxpowerdn : in     vl_logic;
        digitalreset    : in     vl_logic;
        dispval         : in     vl_logic_vector;
        dividerpowerdn  : in     vl_logic;
        dpriodisable    : in     vl_logic;
        dprioin         : in     vl_logic_vector;
        enrevparallellpbk: in     vl_logic;
        forcedispcompliance: in     vl_logic;
        forcedisp       : in     vl_logic_vector;
        forceelecidle   : in     vl_logic;
        invpol          : in     vl_logic;
        obpowerdn       : in     vl_logic;
        phfiforddisable : in     vl_logic;
        phfiforeset     : in     vl_logic;
        phfifowrenable  : in     vl_logic;
        phfifox4bytesel : in     vl_logic;
        phfifox4rdclk   : in     vl_logic;
        phfifox4rdenable: in     vl_logic;
        phfifox4wrenable: in     vl_logic;
        phfifox8bytesel : in     vl_logic;
        phfifox8rdclk   : in     vl_logic;
        phfifox8rdenable: in     vl_logic;
        phfifox8wrenable: in     vl_logic;
        pipestatetransdone: in     vl_logic;
        pllfastclk      : in     vl_logic_vector(1 downto 0);
        powerdn         : in     vl_logic_vector(1 downto 0);
        quadreset       : in     vl_logic;
        refclk          : in     vl_logic;
        revserialfdbk   : in     vl_logic;
        revparallelfdbk : in     vl_logic_vector(19 downto 0);
        termvoltage     : in     vl_logic_vector(1 downto 0);
        vcobypassin     : in     vl_logic;
        xgmctrl         : in     vl_logic;
        xgmdatain       : in     vl_logic_vector(7 downto 0);
        clkout          : out    vl_logic;
        dataout         : out    vl_logic;
        dprioout        : out    vl_logic_vector;
        parallelfdbkout : out    vl_logic_vector(19 downto 0);
        phfifooverflow  : out    vl_logic;
        phfifounderflow : out    vl_logic;
        phfifobyteselout: out    vl_logic;
        phfifordclkout  : out    vl_logic;
        phfifordenableout: out    vl_logic;
        phfifowrenableout: out    vl_logic;
        pipepowerdownout: out    vl_logic_vector(1 downto 0);
        pipepowerstateout: out    vl_logic_vector(3 downto 0);
        rdenablesync    : out    vl_logic;
        refclkout       : out    vl_logic;
        rxdetectvalidout: out    vl_logic;
        rxfoundout      : out    vl_logic_vector(1 downto 0);
        serialfdbkout   : out    vl_logic;
        xgmctrlenable   : out    vl_logic;
        xgmdataout      : out    vl_logic_vector(7 downto 0)
    );
end stratixiigx_hssi_transmitter;
