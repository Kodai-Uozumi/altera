library verilog;
use verilog.vl_types.all;
entity arriagx_hssi_receiver is
    generic(
        adaptive_equalization_mode: string  := "none";
        align_loss_sync_error_num: integer := 4;
        align_ordered_set_based: string  := "false";
        align_pattern   : string  := "0101111100";
        align_pattern_length: integer := 10;
        align_to_deskew_pattern_pos_disp_only: string  := "false";
        allow_align_polarity_inversion: string  := "false";
        allow_pipe_polarity_inversion: string  := "false";
        allow_serial_loopback: string  := "false";
        bandwidth_mode  : integer := 0;
        bit_slip_enable : string  := "false";
        byte_order_pad_pattern: string  := "0101111100";
        byte_order_pattern: string  := "0101111100";
        byte_ordering_mode: string  := "none";
        channel_number  : integer := 0;
        channel_bonding : string  := "none";
        channel_width   : integer := 10;
        clk1_mux_select : string  := "recvd_clk";
        clk2_mux_select : string  := "recvd_clk";
        cru_clock_select: integer := 0;
        cru_divide_by   : integer := 1;
        cru_multiply_by : integer := 10;
        cru_pre_divide_by: integer := 1;
        cruclk0_period  : integer := 10000;
        cruclk1_period  : integer := 10000;
        cruclk2_period  : integer := 10000;
        cruclk3_period  : integer := 10000;
        cruclk4_period  : integer := 10000;
        cruclk5_period  : integer := 10000;
        cruclk6_period  : integer := 10000;
        cruclk7_period  : integer := 10000;
        datapath_protocol: string  := "basic";
        dec_8b_10b_compatibility_mode: string  := "true";
        dec_8b_10b_mode : string  := "none";
        deskew_pattern  : string  := "1100111100";
        disable_auto_idle_insertion: string  := "false";
        disable_ph_low_latency_mode: string  := "false";
        disable_running_disp_in_word_align: string  := "false";
        disallow_kchar_after_pattern_ordered_set: string  := "false";
        dprio_mode      : string  := "none";
        enable_bit_reversal: string  := "false";
        enable_byte_order_control_sig: string  := "false";
        enable_dc_coupling: string  := "false";
        enable_deep_align: string  := "false";
        enable_deep_align_byte_swap: string  := "false";
        enable_lock_to_data_sig: string  := "false";
        enable_lock_to_refclk_sig: string  := "true";
        enable_self_test_mode: string  := "false";
        enable_true_complement_match_in_word_align: string  := "true";
        eq_adapt_seq_control: integer := 0;
        eq_max_gradient_control: integer := 0;
        equalizer_ctrl_a: integer := 0;
        equalizer_ctrl_b: integer := 0;
        equalizer_ctrl_c: integer := 0;
        equalizer_ctrl_d: integer := 0;
        equalizer_ctrl_v: integer := 0;
        equalizer_dc_gain: integer := 0;
        force_freq_det_high: string  := "false";
        force_freq_det_low: string  := "false";
        force_signal_detect: string  := "false";
        force_signal_detect_dig: string  := "false";
        ignore_lock_detect: string  := "false";
        infiniband_invalid_code: integer := 0;
        insert_pad_on_underflow: string  := "false";
        num_align_code_groups_in_ordered_set: integer := 1;
        num_align_cons_good_data: integer := 3;
        num_align_cons_pat: integer := 4;
        phystatus_reset_toggle: string  := "false";
        ppmselect       : integer := 20;
        prbs_all_one_detect: string  := "false";
        rate_match_almost_empty_threshold: integer := 11;
        rate_match_almost_full_threshold: integer := 13;
        rate_match_back_to_back: string  := "false";
        rate_match_fifo_mode: string  := "none";
        rate_match_ordered_set_based: string  := "false";
        rate_match_pattern_size: integer := 10;
        rate_match_pattern1: string  := "00000000000010111100";
        rate_match_pattern2: string  := "00000000000010111100";
        rate_match_skip_set_based: string  := "false";
        rd_clk_mux_select: string  := "int_clk";
        recovered_clk_mux_select: string  := "recvd_clk";
        reset_clock_output_during_digital_reset: string  := "false";
        run_length      : integer := 200;
        run_length_enable: string  := "false";
        rx_detect_bypass: string  := "false";
        self_test_mode  : string  := "incremental";
        send_direct_reverse_serial_loopback: string  := "false";
        signal_detect_threshold: integer := 0;
        termination     : string  := "OCT_100_OHMS";
        use_align_state_machine: string  := "false";
        use_deserializer_double_data_mode: string  := "false";
        use_deskew_fifo : string  := "false";
        use_double_data_mode: string  := "false";
        use_parallel_loopback: string  := "false";
        use_rate_match_pattern1_only: string  := "false";
        use_rising_edge_triggered_pattern_align: string  := "false";
        common_mode     : string  := "0.9V";
        loop_filter_resistor_control: integer := 0;
        loop_filter_ripple_capacitor_control: integer := 0;
        pd_mode_charge_pump_current_control: integer := 0;
        signal_detect_hysteresis_enabled: string  := "false";
        single_detect_hysteresis_enabled: string  := "false";
        use_termvoltage_signal: string  := "true";
        vco_range       : string  := "high";
        sim_offset_cycle_count: integer := 10;
        protocol_hint   : string  := "basic";
        dprio_config_mode: integer := 0;
        dprio_width     : integer := 200;
        allow_vco_bypass: string  := "false";
        charge_pump_current_control: integer := 0;
        up_dn_mismatch_control: integer := 0;
        charge_pump_test_enable: string  := "false";
        charge_pump_current_test_control_pos: string  := "false";
        charge_pump_tristate_enable: string  := "false";
        low_speed_test_select: integer := 0;
        cru_clk_sel_during_vco_bypass: string  := "refclk1";
        test_bus_sel    : integer := 0;
        enable_phfifo_bypass: string  := "false";
        sim_rxpll_clkout_phase_shift: integer := 0;
        sim_rxpll_clkout_latency: integer := 0
    );
    port(
        a1a2size        : in     vl_logic;
        adcepowerdn     : in     vl_logic;
        adcereset       : in     vl_logic;
        alignstatus     : in     vl_logic;
        alignstatussync : in     vl_logic;
        analogreset     : in     vl_logic;
        bitslip         : in     vl_logic;
        coreclk         : in     vl_logic;
        cruclk          : in     vl_logic_vector(8 downto 0);
        crupowerdn      : in     vl_logic;
        crureset        : in     vl_logic;
        datain          : in     vl_logic;
        digitalreset    : in     vl_logic;
        disablefifordin : in     vl_logic;
        disablefifowrin : in     vl_logic;
        dpriodisable    : in     vl_logic;
        dprioin         : in     vl_logic_vector;
        enabledeskew    : in     vl_logic;
        enabyteord      : in     vl_logic;
        enapatternalign : in     vl_logic;
        fifordin        : in     vl_logic;
        fiforesetrd     : in     vl_logic;
        ibpowerdn       : in     vl_logic;
        invpol          : in     vl_logic;
        localrefclk     : in     vl_logic;
        locktodata      : in     vl_logic;
        locktorefclk    : in     vl_logic;
        masterclk       : in     vl_logic;
        parallelfdbk    : in     vl_logic_vector(19 downto 0);
        phfifordenable  : in     vl_logic;
        phfiforeset     : in     vl_logic;
        phfifowrdisable : in     vl_logic;
        phfifox4bytesel : in     vl_logic;
        phfifox4rdenable: in     vl_logic;
        phfifox4wrclk   : in     vl_logic;
        phfifox4wrenable: in     vl_logic;
        phfifox8bytesel : in     vl_logic;
        phfifox8rdenable: in     vl_logic;
        phfifox8wrclk   : in     vl_logic;
        phfifox8wrenable: in     vl_logic;
        pipe8b10binvpolarity: in     vl_logic;
        pipepowerdown   : in     vl_logic_vector(1 downto 0);
        pipepowerstate  : in     vl_logic_vector(3 downto 0);
        quadreset       : in     vl_logic;
        refclk          : in     vl_logic;
        revbitorderwa   : in     vl_logic;
        revbyteorderwa  : in     vl_logic;
        rmfifordena     : in     vl_logic;
        rmfiforeset     : in     vl_logic;
        rmfifowrena     : in     vl_logic;
        rxdetectvalid   : in     vl_logic;
        rxfound         : in     vl_logic_vector(1 downto 0);
        serialfdbk      : in     vl_logic;
        seriallpbken    : in     vl_logic;
        termvoltage     : in     vl_logic_vector(2 downto 0);
        testsel         : in     vl_logic_vector(3 downto 0);
        xgmctrlin       : in     vl_logic;
        xgmdatain       : in     vl_logic_vector(7 downto 0);
        a1a2sizeout     : out    vl_logic_vector;
        a1detect        : out    vl_logic_vector;
        a2detect        : out    vl_logic_vector;
        adetectdeskew   : out    vl_logic;
        alignstatussyncout: out    vl_logic;
        analogtestbus   : out    vl_logic_vector(7 downto 0);
        bistdone        : out    vl_logic;
        bisterr         : out    vl_logic;
        byteorderalignstatus: out    vl_logic;
        clkout          : out    vl_logic;
        cmudivclkout    : out    vl_logic;
        ctrldetect      : out    vl_logic_vector;
        dataout         : out    vl_logic_vector;
        dataoutfull     : out    vl_logic_vector(63 downto 0);
        disablefifordout: out    vl_logic;
        disablefifowrout: out    vl_logic;
        disperr         : out    vl_logic_vector;
        dprioout        : out    vl_logic_vector;
        errdetect       : out    vl_logic_vector;
        fifordout       : out    vl_logic;
        freqlock        : out    vl_logic;
        k1detect        : out    vl_logic_vector;
        k2detect        : out    vl_logic_vector(1 downto 0);
        patterndetect   : out    vl_logic_vector;
        phaselockloss   : out    vl_logic;
        phfifobyteselout: out    vl_logic;
        phfifooverflow  : out    vl_logic;
        phfifordenableout: out    vl_logic;
        phfifounderflow : out    vl_logic;
        phfifowrclkout  : out    vl_logic;
        phfifowrenableout: out    vl_logic;
        pipebufferstat  : out    vl_logic_vector(3 downto 0);
        pipedatavalid   : out    vl_logic;
        pipeelecidle    : out    vl_logic;
        pipephydonestatus: out    vl_logic;
        pipestatus      : out    vl_logic_vector(2 downto 0);
        pipestatetransdoneout: out    vl_logic;
        rdalign         : out    vl_logic;
        recovclkout     : out    vl_logic;
        revparallelfdbkdata: out    vl_logic_vector(19 downto 0);
        revserialfdbkout: out    vl_logic;
        rlv             : out    vl_logic;
        rmfifoalmostempty: out    vl_logic;
        rmfifoalmostfull: out    vl_logic;
        rmfifodatadeleted: out    vl_logic_vector;
        rmfifodatainserted: out    vl_logic_vector;
        rmfifoempty     : out    vl_logic;
        rmfifofull      : out    vl_logic;
        runningdisp     : out    vl_logic_vector;
        signaldetect    : out    vl_logic;
        syncstatus      : out    vl_logic_vector;
        syncstatusdeskew: out    vl_logic;
        xgmctrldet      : out    vl_logic;
        xgmdataout      : out    vl_logic_vector(7 downto 0);
        xgmdatavalid    : out    vl_logic;
        xgmrunningdisp  : out    vl_logic
    );
end arriagx_hssi_receiver;
