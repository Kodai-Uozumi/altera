��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���a?K���J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-~09h�i�Nq�{5��]�0�lK'���Xw����Q4f����om2�YQ}�U�"g%�\�Ji��'��%�a�z�o���Ή�����f�p��G�42c�Ϡ\�)zL͊�q�� �^�ߏ'ER���c&;\e�L���'��-d�Ry��\�v���T�©ޒ�����s�VKOi�~�n�
���b����Y�{'%s4C>-��3v#��.X���*"v%)�����iR˳͠m�xW�g]����n(���˧[(X�#��§S6]Z���榡dB� L�s;X�a\�/���~09h�i�Nq�{5��]�0�lK'���Xw����Q4?���ʢS����E@�gh1���Yh�\��q,f$�7Q0- ��Ck�4���_z�k�۸�y�uZoO�=���t8� L�s;X�N�N���aC�h�>��!�̰���_8\/HiO���L�~h0%�������E3u�;5B5Y+��q	k���A�XWf^64W��^�o�A���,r�s��pK�����o���M��JVLM∓/^
wUgJ��Kʸϸ�N�
�o��djf[P�O�+`�W��� ѦV��7^�9 �;���b��iAj %�Ho�-[�v:v�o���+����7X��U�?	r���g�0�u�w��$C��׫�J�є^ֻ����XP���-O/ [р$	3�Ð�9�X�e�b��@�zL͊�q�����芶t���6��^hq��:�y���OJHn��z��r9�3ꓩ�l;��!I/�������A��1��+�W�Ń�I��-Ndp��5MYu��>��
��������0��8���o�5���ڲ$ Zh0%���ԛk%��q{�f��a�t�v�5��m��K���x�k�@�1z�:맷�خı�)tp8��x��ƍ���<$��Q��[�y�3�Y�`�'n�^0oW��T^�<��Ƶ�L�9����#i/G$[�����b�QO�!]���pxq{�f��a�P9b�� ����X�[$��Q���N��T����b�QOu��
Q��x�$<���GzL͊�q��[���0e��㎟�>z�����r���E�sy����.G�}���fŧ���|���x��EP��\|��EaV�5�j��l2�bczL͊�q�� Ky��:~�)1:���iR�@>���:����{��Ƀ��-jD^�o���"�PЭ��i����Z9p�����1F�mq{�f��a�6T{��2~*.�P[k�KW�*�	S~�i25��[%��4�[ⱸ�ND[�Q0��U-^G���c���%���+��q��N��^,�p/�����c�9�:&�ߦ8���Hm�č�Y���S�)37J*uV��4�����k�b���9/���`���6j����ƛӧ�#2�|���˿x�"�,�>E��<��z��}���<���_j�<)G�9� ���jZƇ$�g��U-�eHe.S:�w)��=�sEټ�O
�_�Z)���Øf���Q�0�	�����T���9�dMbZ鎬����)pq��Hj}��0>�%��WT�j
�I��w��,c�A�L' &�M���=�sEټ�*��T�����`y����Q�C^��z�s[e�t��`�0�דPg�'|����d�k�(+\�(_7MԲ�����{l�f|����%Hlܼ��2��}n	�Z^�t���,2����X�kX������`4�E%v�~������]�!�����#e���5��(_]�Jg����-c �ЄW:'�|�9+R��2$6�sIw!
�h9RE]1L�D�W�D�b�v�~������]�!�����#e��_:�Z���,2�����^���@�d�_C�VJ����̕���(��h�9�@��p�Ia��ܛ8�7�FG<�`�hE���Mz��;��ҋX����0�a1i~Js9}B�Ź��ݏ1��𠛕!��L�ވ���ۭNJ?�s�C�,������[GL�����K+I�\�q��N��f�;�>)�~�`�0��|��].��'���XwSg0�#�aea���||��/8'�G~+�3;��\���\��k�zph5)�� �;7mg�o2��c=�_R�k��������ǈݻ�:������<��z��}�צ:�)1q7{�q�B*�2���u���d���=A�2�S|���f?��� <�"��=aet�V܉i��d�=i"}�۞h�G��+^zO��!n}y���q���U�J��ZvA� ���ѡ�e�LZ\^�e���Eы�`�M7Э���j��S��^1�)��ܘ�b2��c=�_R�k�������I�}j����CX�ҋX����0�a1i~J�!������ݏ1��𠛕!��L�ވ���ۭNJ?�s�C�,����&�2 ���������x��lV��(C6	�YI܁���!n}y���q���U�һ�aRp�� ���ѡ�e�LZ\^�e���Eы�`�M7ЭH$#5b ���Z�s9�*�@w�[�u=�@X�wZ K�Ϋ�v�~������]�!�����#e��,�SVj]�Jg����-c �ЄW:l�mq���)�:V�7	|[��
ҦV�	�o�Jr�)L�/��Ĉ=�t��Hܯͬ8�.��č�Y���S�)37J*uc�A�L'�f?S��|�b�@a(􆿳�ʨ�6�j���L�9�r.p�B*�2���u���d�ӿ�>��f]��A�5�D��o�Pc��?@W��o�BѰ_�Du\��-���(���5������:�TD���rs�i��=29��a\e�L����owђN�~��&�t�).?-��o@�e6qR5L�/8'�L
�2�Ot����F�2�v����o/�;�����=f��9c����3���S�����E#񲇽t8k>6s����]�!��R?��bgR8�Ņ�~L�e�LZ\^ �@'�ZX8�5}7�4�B��ٴ%+����#����ir�� �:&��k�t���.鶇�?6� ��|7�>P�2-i_���F���-����gۏ�#��:V^����9�%a�E�IO�2_�ⷱ�ْl��]�B9�θ�c}k5�Y���[}\w��B���Y��]����MT�	��y���!�`�(i3��W0i��^_0;%]a}�� �с�$��R�lD�"5� �S�jn�Ł�K紣�	��h5����Z�>)��oz��KUq���8�/>�"�Ax=]A��O�T�`�[����)=��%1�{�C���g#B��F�!�`�(i3x�]�V��\#O���oӧu��՘�uw�@.�/wc1����#�F�!�`�(i3�o��C!T*Y�{'%sJ��m���P�)��j����16X��5@~Ju9gUS��������[�=9t*�e+��4<��z��}�<ͧ�:|f;[����"���.��E����F�ҋX����L$�����/'٥��gV؞� %�0Y%T��BPS�)37J*uc�A�L'M�;��p�A��.�'f3�T�\ ���YP�UZ���*l�86Yl���#�]�!��	Ǹ�y85�V��t����.&H\�HP@�a����U�p��
���)�"���R��� VU+I��(�@$.>��K����\#+��Sз��x��@���U@���:��F�ʳ�A~�0 �i7�sp>4��D��6ʜ耚ҵԼ�\�v�)��+�}��l���n�2 �.��c��\�vŒO�����i#@���%&E����T�OL�Wr��k��&�8�ҋX������S8���<ށ���h���o�8���/����42	vX�7P��T�<��z��}�Q2�+�Y�r���}�č�Y���S�)37J*u)T{6T'�n�<���v�~������]�!��V�,�q^����Ho�d��!n}y���q���U����7Y،���Ig`i�ҋX����@�ڗe'ٜ�U�n~q_3#ڸZ鎬�����c[��/n��9�n��(�
t�������2����U�p��
���)�b���"v����Ɛ�,�)�H"�Lܛ�ð��D-�]|�8M͌4s+�nyz��:W_Jܛ�	��|��	(���zL͊�q����#N��#^�Vn1�*_��h��~|K6�[T�)���}0�st&���\�v���T�©�'�3�$ �#^�Vn1�*_��hзܽG��?2^�9<o�nïi�JHn��z��k"����_i��Rp�������О.[<՝4��&ˣb�O��'F,�����r�|S���?˻D?a�G���6(:�*4�?�^ֻ����XP����� ��p�FQiҗ�.���t8��U]�lEGV`28��4xc�\^��d4\��N(�RZ(�󕏜9��㮑�ToE�(J�qE^q{�f��a��4�6�tږV�x)"-��齚ϦM=�S_!�:d�=�k2B]p�"m���C�,���3�.JHn��z���T��Ćm���n�ٟ��f��#����bs�������]��5��f�4
�Ǽ
Ձ����&��_�G��GJHn��z�_c)���8��%�a��/=�c ��%
��(T��5��8�t��\�v�CF���y7�5����`Kx���T�LEY��]-� T2��zL͊�q��e�[,E�Ћ�l�TQo�RGw�փZ���0�JHn��z���z�O҈͌4s+�nyg__{���@O
�`z0�KP�i�IÙ=�H��K�)�PMI�������@
/���%
��(TyT��V��Q`��J��k�=[�p�����.�q�-���Zxq��:gB(q�'T�� �������?˻D?N6ߠ������?!�KW?���#\rgd�TpubMpIÙ=�H���n�����U���%�G�܃?���1#�i�0�o�݀�̆����E��nU\T�7Z�#���b����8�MN)�j��&!��"�F������mj�pzl��a�� �܈~\�Mf���9���q���U�?�����"2�#�>��~���1��B����qC�<��1���?��;���H��Ig`iZ鎬�����7]=k���1�&"i�9�����>l\�}�jT%q�#��]�!���äs_���l�mq��L��T��>�]bU9]M(��۷�_,2��K�QY/����[B�����'���Xw�P>a�.����'�#&�3��3�-��y��hi=O��s��#%��$�z��e�K���d�٣���-��� ��d�_C�V��pµ�Ս��������K+I�\z�f�a��c�������7P��T��]�!���äs_���l�mq��L��T��>��Nv|��U+�ei�Dj�������8k��t�7P��T��]�!���äs_���l�mq��L��T��>���VuS!ִei�N�iP+�����u�	NMf���9���q���U�?�����"2�#�?�< TL�MT�5B�������;Q�U	t��c��`ʗ�Mf���9���q���U�?�����"2�#�?�< TL�M�����0� :�]4�W�{Њ�l�L���9M[B�����'���Xw�P>a�.����'�#&�3��3�尡�������;Q�U	t��w��n��y[B�����'���Xw�P>a�.����'�#&�3��3���<�4������;Q�U	t��\�T~�SMf���9���q���U�?�����"2�#�?�< TL�MK}�V�h�;����;Y�hg�N��M���5^s��Z�-��ݾNt�Yӑ!�;�?��R��V�
�]�$��'���Xwa'�<� \�_Q路�9�ͤ3�G�ҏZ���]�!���1����mӑ!�;�?݁*=���$Ak6�r),�d�٣���$�j��ш7�����R<�#)��Ľ=
Q�¸�)�`E5U���c@��`Xg?�����Y�Y�{'%sgeߪ�{��EA��*��ʄ6�PǨ�o*� 7�v�ԯ�o��f��)�`E5U���c@:��!�6�F���D����'���Xw�j�7��x���T�X~0���2Bm��Z��,0=]^	�&QR�u9�����K�Q/8��A0��Ig`iZ鎬�������(���@��/��
x�GM�
 /R�1屖ʨg��U-�e9��K哧-�
�W^޺���!� E�����Z鎬�������(���@��/��
ђ{)8A�^�V]��}%鯅�pzl��a�H/�I��!#��L�$E�����'���Xw�j�7�����n����H�HoLf,0=]^	�&QR�u9���G ��7O��E�&����f��jvr��Q������h����@$˺/t��꫕qŧo��K�O`�Y��
eU���c@cy�@�Xŕb!��u�PQ�>\Ճ�<^	a
$����$�Q�r �K��Im7��JL���Z'?��Ǌm����0�E>Sx�lޞ�ό���.���K�Q9�ͤ3�8�iE����P
Z鎬������Ȥ�8��P	X���������7��s�KTkѶ���� �Cs�9`H�玨��Sx�lޞ�ό���.���K�Qbs4�U�y��z��~�՘�=Y��_�0z�cUL�����t�kI+a����R�1屖ʨg��U-�e(�!W�4���*!��Uk�e~���G��[�֔�	�_t�����j�u���
�����ﻋ-�����S8��J���o��Wq�;5̠�&A���T�\ ���|.�Tӏ:�L�
�+��[��XMf���9��Y�{'%s43u�R��V^[s-�H��4��j��
�ߴm���&�t�)ɝ:���vvN�c�������ᖚQs��m6�eIOkѶ���� N�B.D��z��a7��ﻋ-��ȳ�Ǿ�����"y����7�)=�lv7�H^%o�Z��beNY� o����[�c�Ĭ	Mf���9���q���U����ۑL��YL�P���-w˕���?����a�x��3����Hhqu!���5�Nn���4L"�#W��xW�Kg!�h�����7�$�G�j/����X�e�zP����=���m\Ӓ�qܛ�	��e�N��W�M��0�d�Sd��_�a���n�|W4S�8Mi�K�z;�"�nT��z��uWU4y5=>F/ġ"���Չ-d��r�b+ӄ�bİ��i+��*�I�GIN�|L9_~��O3m�M�n����x5=��{t_�sVh�a�ohWt�_a�1�܄:h	}4���!�fJ��l߮�pd�Zз���?̕U�/j�g4A���{0Yafk��r.y����nL���~C�V�T��a׈Eg#f�z�q���<�{�!���"�ֱ��R8v��j.Z��$�sӢ�]3�����c��(r$����Gd"��U"�̩��k&Q��8�'��j^ҩ#��u1&2�%�	[2�����Vc2�����Vc��Y7�z�p���w�nrm؊(�p��Aby�2�����Vc2�����Vc���1� -N&ݨ)�����a��	{��#-�	=��>QH[[����q�f��6&1�1�<Y�W�q]=`爼#��8h� 1�����f�c��k�-����B���f�;�>)�(���Yr�r��`�^�qFQXI�DZܤ�jh"r��RǷe�b��1j�L�uVBդ(m�캧xӍ.��L-�yC³RǷe�b��1j�L�uVBC�9mE_ݧ�f�;�>)�M�?��?+�r��`����s7b`?�'n��c�,�[`�t���iqFEĈ�d�1r6y_s� ��DZܤ�jh"r��c,W� K91j�L�uVB1��0�캧xӍ.��L-�yC³c,W� K91j�L�uVB+�o'���<���I�&�`E�b�.�.oA!�?2��l��Y�Q+�zN����9�2�L�1�,I�v��e}0�E�g�������(ӈ��\#@��\2�����Vc2�����Vc2�����VcREBR�hHr��쁳.ۤ�a��:[\�����
�N�1�� ��2�����Vc2�����Vc��`���4>V~ya̋o�C�!�2]�oک�C,@���w��XS9T�c}���W>ܛ�tU��.���D�k��5L1膒��5��R
2?a)���*=���$�����-?2]�oڄ�7amL�#��M}��R��	π2�����Vc�cRq>h���迴ކ��	uz�t��f��I�2�����Vc2�����Vc؁�Pu�5���<������+�o�T�a_�wj��\f��x��±eKr�V�f�tށ�W����`�n��U%aWp��.�替��+���<j�2ʧ6�0�h	��6�y/�
x���0�o5�����EO�{����F��l�}��=�sEټ�K�2��M�
+,I�2Sj�	�$ɜ����0+C�%�_�UK%=k�Rm����?�I���6\�4�@���(�?<-M�O��~��i��"u��Y�H�-z���t˨{��-�C��7u#md��9�ͤ3�8���~կ�@/��r �)������I�ɔ)�([��}qn
V~$�V(�z%^�F�_	*��݄���8�Xr��?��Ǌm'r�_�(p�Z!h�-'�X~0���2Bm��Z��,0=]^	�&����ג���a�z6�ZǢRMlC�b~*��s�ai^w&����|-�se�Pع���a�	�+4D@��9�Uz?��Ǌm'r�_�(p.�Sx@5Mp�s��L����qM�&����1���n��	�d��-��!rϚ���Z�B F-W�����@/��r ��JR��W�xU���c@:��!�6�F��h�G��W?��Ǌm'r�_�(pK���L���4�04�jfx(�i��/Rh�x#�L_�(D{ͬ�y�4����K�K}�$� ����T�H/�I���x~bCu����
wcҴ�x�#���c|B��y^X,0=]^	�&QR�u9��⍬�|?�O	�#�O�l�1C��(�H/�I���΁�4���p�ɟ�Vk2�aI��[�n�g3��9�2�L/8��A0�/������kkdBө�3�*{�����<��ї�^ˑJ�|\�
�?ќ�jw�jV��WD�@��/��
� �j<�Re�Ŵ#����#g�k��g?	��oc�Y�y9�ʝ�)H���g�0�u�UӇ�_�,����,|up�LXS�˷��{H�3)-7�ٙ|p�� ,�;Rt���H�.���\+q�+0�u�fF�5.]��۪	�}a4����@[�_zβrrZ�0m�\��A�.4��M�H��px�]�5����V�X~)v�0����2F�����b�QO�
G<�K�!�T�.���gڟ4�{"�Lެ�kJ�9#���ޕ���6vD�Λ�{��x�l��1i�t�U0_�=2�?�.��}@",|up�LXS$�؁�QG�%<��>�@V�� ��n��i�a�\��@�n��Wrȿ.\5�Y���[}�r�U��vL<��x��±eK��K�x۶�*U*�������S,�D�c��Q�e�ȵ-O��l�@jen���F W��!��r�l ����xl�@jen�-���<86ꕅ|ںi�����s&���EO��J$H/�I��]�=��&\�8qTmI(x;��|B������X~)v�0���"�$��'�Hm��1�C�G���-�����؍R?�6��'�|,kW�A��ˮ��V�rsSRąf�c~���[1�
�8jYj���W*�C��-^��������>��E�V�*Oб�ne/���d}��[�ƭM@m�gwg͇�WDv�b��'�s�ɧ�E�\'��fHXz�'�z?XÚ
�3]Pm��KCw.���>��gO�����h�ZnEw�S��EC��Us�_��s�֙�M�˵·|���d� ������TU���c@�鼱�v(h6j�"Hs|aqV���[ⱸ�ND[M:b����`.��g�a0��I�l����)�u��ݵdw3{���yu��mDrv�<�2�Ҧ1���Z�וzj7i�j�ʜ/�;�o1[��wEGͶ0h�5e��`'��<��Ȝx��y����ү�+ҋ�y�$:����!� o[v<�FH/�I��t+�FQ�X�J�1���۪	�}a4������s���5�`_�ʵ�1BJ+�Z���"5��������Q@[�_zβrZ�tH�=���.�˕1��@���j����T�OÈ���)�l*ªK����'�(j`N���Ew�S�����p*)�*C�8؉b�'��(�~��e�.5�����O2��_E`s��E��"���h�=���������!Z�*_#a�u�CRXp-y#��埄��)�� G�/~ޖ+�x%��ό�;�LȫԷ�/����t��2�����Vc2�����Vcl��w&� 1ᗟ��ÝO.ZR=���<� �z9�GKP�2�����Vc2�����Vc\��H;�21h��ʠU��jyc+j�H/�I���x~bCu��O��/ӎ����L�I#5𵪋��S�%�i��:�}��E5�%��
~�.as�Y{h����Y'��y��f8�p!!k�^/�&@�d��w��������\Y��K�,h��j�3���v`�%����5/:�� ��N[��ڇ�8�@�mh@�!݄�j}����f8�p!!k]�<����K�#ln3�ɬc��WN��gE��ң]=��j�F���+�= �i�,Z	�FWJ�)T�����������6<k�r�Q�#�ix:���t��9C����#;�ec��Uioέ���'*$�T���@yx��)�� G�/ސE}yޱ;��|B* ^���x��obV��|���d� ��Z<��C�f8�p!!krD�؃���L�C���ea�Xi��T���H�*h����L8�&a;��|�v ),�?���#�R	[����Kv� �~�9rF`_�ʵ߶��57�'�[b%Ɨ��������!���?t��my$�N���4H���rw�&�z<a��N� φ��<�6�Ps_*�GqW�w��fD!��I\+������BL�R�pM���#9Wٓ�6��<��7��qib-)\����]���#9Wٓ���2F���\|��EaV�5�j����x`u�P_g3���K����'�kk~�AD���Z�וzj7i�j�@���-�qx�'|�9��x~l��Uh����L8�C�	R�x�������ՙ�.�h͉��7,F��[WL��g8!�|!��[�N�g�c�`�zc՝Rq��R�ҾGmdN�<@Iv����-�T�8��e�[b%Ɨ��������n�+7���ߦ�����q��>^��x(�i��/R�*�W�Ǹ!2�͞nOY�c�����t��7Y34뙩A��n�4�uVYY����!�͒C@�~TĪj`g���5���%���1�_G �1w�{�kH�K���,"b��j�3���;n�c�S�S�W1�9���ᢳ/z��I5�	�����AC�	&}w|�"��P�9��o�1��~��\o���x�
�f��Yu�]bu̎,+$\�M�\��}�NQC�U�y�`D}��I�fQ7�H�8i�H�玨���$���:�%���2F���\|��EaV�5�jr��X�^88u�P_g3���K����'�Ŵ#����#g�k��g?	��o/�#��J�d�{��8Bl $���n?3NϜx;��c�� N��r*�Ɠ�d�w��$��*of����Kͽ<\��-M�O��~��E��5���VLpW��I+a����R�1屖ʨg��U-�e�:>r9�*v�ߦ������Z?�>0=�Q`��J��G\O�E朦����Uh1�-���)+@����(�8#�H��71ri���ђ{)8A�^�V]��}�dh_��tCdN�<@Iv����-�T�8��e׏�����MFi��|ր���5V��	��yo��Rn��$���\�uB�3DO�9�?B01�|2 �F�m�+2G\�j��fxŪ5eOt'ʽe��jV��WD�H$[4D����ɣ��سH�O�PWy��g�:2�W�(F���E�,(W�;��|B* ^���x��obV��|���d� ��Z<��C�f8�p!!krD�؃���L�C���ea�Xi��T���H�*h����L8�&a;��|�v ),�?���#�R	[����Kv�<)G�9� �H�HoLf,0=]^	�&��[�4�f,�{_8�Y�����t����-���)+@����(�8#�H��71ri���ђ{)8A�^�V]��}�dh_��tC�E�VmM���d�{��8B�<)G�9� �H�HoLf,0=]^	�&����ג�J�1���۪	�}a4����@[�_zβrꢯ�wv��\�j��fxŪ5eOt'ʽe���F���✁���l5v�I�DSV��JM;��s;�Z����(t�	H�޹q��}����M)�*C�8؉b�'��(�~��e�.5�����O2��_E`s��Sf�%�����.i$ۇ��;"�1���dUl��3c��)��HS�kGQ��s��9P/1q���<�{�!���"����F��2�����Vc2�����Vc2�����Vcl��w&� ����e�<9�ǆ�K�<^&!!HY��f��I�2�����Vc2�����Vc2�����Vc��%3$��|�-@2����؄V��^��,԰^��:S	m���cbp��'@
9��y�uP����.(�g���N�\[�?�����l����4�n���xǊ�6P6x]G�H�޹q�ֶ��}�Y�j���@+�b���-~�*���t_!0h��(Z+�<Vo�eo0C��:�4�*��2�hil�C��3�I2E�D�����&���V��h4����O�$��do�����z���R�V�x�;��l����4�n���xǊ�<)G�9� չ|Jo��Rx���T�LEY��]-��b�;���Y�d�X���l����4�n���xǊ�<)G�9� U�G�@m<��WP��F���q�2�	%}RN�y]I�Eۇ�m���5���7�#�x�-��:�.�zΑ��$��N��E�EX̦,\ަ�It*���1��ͫ��;���^hq��:�V��ÑR ����*��Y~��`�J�(��Q|3�'�2%$>�	}o2���Q����$0��b�;1?�[F�sp֟kh��b��	���U(���R�X��Uq2��Z^��:8�~[㧼������L��S-���"h#�)��!��ZB�;�H���o(�,ebY�s�3|�&�Z�oO�q��rH��i�׻�Z\�i�æW���h�R�⿣:�d���φc�����7Y،��!��ZBϵ��=%1v����ƾ+r����%< ͗���{�T���^A��3c/��!S�!��LBٜ�U�n~qbS�xǠ�jP"F0�4�fn��9�nD�m	$��\Ef�>:��;���Q>�^2�����Vc2�����Vc2�����Vcl��w&� ��tF��J�����{��ܨ���[����9�GKP�2�����Vc2�����Vc2�����VcSd�*-}Q�O���ƻoW��	]�	�g��>���,���Ks�=E��r�Ø}[�S�>=k�Rm���<��=����7�j�Γ�N�g�c�`w��J���m���=+�"ª���#Â��&?�i#�z h6���{���I�q����.Z�2{4x{^4��*m�D�$0��wO��N�@/��r ��JR��W�x�&�jW� ��|�5���+Z�J�1����ݾ-/�uu��ڿ׏�����M��ܐ�}��t�l���Lq�"��2�L������W�p��S,�a�r�ǯ3�4������_ 	>��M���5^s���@�Ę��!{6�R��V���u�g/QP�y����b(�=Y5��Y�H�-z���t˨{�'�ɚe�4����0�E>tT$H�;d�^�F�_	*���x`�CϝQ����\Ef�>neb���.�m���=+��A\/i��KX��iko����Ӫ� Q�����([��}qn
V~$�x2�:��N�B.D��o}����ĳ�e��@Q��K,8cU���c@�H��	W��N�g�c�`�4�!���T`��J�^^�F�_	*��[��9���&�(5�;2�f�3�Ұ5ϝQ�����H��	W��N�g�c�`�4�!��䰈C%�>�^=�����o}����ĳT۳�͕���zt��[�A�qL2�cU�:��(�J�1���k_���b_!2�͞nOYգ�-�D��>P�2-i_e����͂�I.��^�