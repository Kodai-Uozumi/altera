library verilog;
use verilog.vl_types.all;
entity apexii_hsdi_transmitter is
    generic(
        channel_width   : integer := 10;
        center_align    : string  := "off"
    );
    port(
        clk0            : in     vl_logic;
        clk1            : in     vl_logic;
        datain          : in     vl_logic_vector(9 downto 0);
        dataout         : out    vl_logic;
        devclrn         : in     vl_logic;
        devpor          : in     vl_logic
    );
end apexii_hsdi_transmitter;
