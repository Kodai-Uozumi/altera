��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���h�k��$�J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-?H)t� �hz2��ƿ� �lJE�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hp���Ť�Mn��X)r����#�L������5N�1 T�V	�tL��	�{�Κ$M�C7y���v6޿���kq����Eֿ�o0��ܧe���5�/���ׇӭ��!�`�(i3[�"5�QJǊö��_��i@�{ۧe[ғr�,�Ōt�}Uٱ�g����.E�^~_|�����{j�G:� ��'��iI+w,A��4�M\���Z ��a�O>*���
��#kz��GN�P�0v���uP!ߌ���^����Wړ��]b�=#;6�#t����nB3�+{Cz��3�<A��d�]��<��&�gG��Hc�e$���=�(v
���O>E$I������T���Q���!i��ӯ�0���&�:�u0&����x2�Zy����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�jM�1}2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!����j.�n�Ax��PR@?�Q|33�����rqn���wѪ	/g�%�W��{�RX�>w�P���u0�������k�V�99^�)�S��uC|Q�����9�ih\���6�oX��s�At�Ӡ�-������u�=�xs�1����";1�(�����]a�{��ۊ�d�k�`�?��<�� ��o�}a�Còz�;^�ru��e��_$߼
�d�YiUbiX>�"��g��3�G��/8'��ި]M�}xf���T��Mߟy�����n��1��\�p��/L�M��Y�Ҁ����r��{��>ڑ/8'�odgƚ�| �����q��5k�^�78���N��ov�Op����	�Y8�>����;% ���W~�_Y�1�����q[��\�jf)�bdZ0o�v�v���O��q�M�4��{i�etWj%h�W�8������8ٓ�j!�`�(i3p]G��>���<�}��x~QTߨ�O3��\�'�y'��BS�z�5&n��ū��@�k�!�`�(i3!�`�(i3!�`�(i3}[x��8��`��Ć?6�!s}6,e �ǟ=EZئ;z&����+�E�r{����JDn ��a�K�.:gdW(o%�)���;t|������D"�~����p�4���='߰����`H��b/3j!�`�(i3!�`�(i3�F{/���!3~�(Z��GmO��%��}�.����M���5^s1@�&'iKb�آ[�~,ΗG\�ʢ�X�=1�����
�^��j"��Q�]f�p����=Qsz����Iv�.�GzEc.������������X�k=o���Fz�!�`�(i3!�`�(i3IB�]�!P���b6p!!v*!���&fB�@��X*,l��d���F6���ׇӭ��!�`�(i3!�`�(i3 lF�Z��f}�y�F�&��S߭;�(6��3{��|o	���=l"�,�>E��&�3�y�2��J�J�T�S1(_�'�&r�~,ptQ��k$Vʴ8X�S����TXP�e�g]�H��֟B��Ўek'`�j�13*�á)ˎ	��[�!%&oA�\ֆ�
'��(�<��
Aʎ^g!�`�(i3!�`�(i3!�`�(i3�|j��"C���ޝsn?V��-Q	�	:����lg\ ����EO�{��ϫ��u�o���q�Z��?��: 0[�T#�l�/Zw������{%hPb��͓T�)��z��z
��K�O�n���^���D�*�Z�J�v$��A�f�y'��BSƹ�#�y�w���	B$�@�A�w{6��(�N��K�O�n8�[ �n�
�CQYb!��uፁ�&�$`8�+DO�n�;4L&�y;U�2y��}���[N�)J��7)�c�0:S��}1yYZ��� ����@	�1i�myh�~�*�.i,����j�Ə���&,���9�tOHn����x���I8I�%-4o��Iu���'�#&��
 {�L<��-�|��e���RB����bb��Ə���&,��+���!XwOHn����x���I8I�%-4o��Iu���'�#&_�:q`��� �Z)}�6!ת���ېư���o���o��V�x�O`BpI�ҽb.j����kѶ���� ���X%��m�Z9a\������0;8�y�%$���r���{��6;)ܟaTo0BpI�ҽb.j����#�2�/D<�L�k��\|�M4��*��J�Y��в}��aC�2V�Vׇӭ��!�`�(i3!�`�(i3I����Ǻ'n;�>�rY
�����+O~%��짐~��.d����"���p|��X^䀸~�W߁�nrm؊(�[���~$�B2���m���-��
�8���?�*���\�Ə���&,Ƿ	DTjE,���6��q@�2��>�b!��u�Z1~�g]�u�+��
~J[����30�A�zc�RhoŜn!�`�(i3!�`�(i3!�`�(i3�M��n���<����lpU�:�ƅf��	��������6��q@�2��>�o����|�sg�2�:��~�^=��D�,<�V�QK�}�9���u����Fz�!�`�(i3!�`�(i3؝�4W���+DO�n��t!I����;R���fǥ�c⠵���طYRdZ0o�v�V#��ب'�����{��6;<� ֭m�_���ȃEE��$(��{�$�˽�Lk�`�?��<��t!I������h+�w��4܆��O�2C��OG;�['*�p!!v*!���O�{�
;����"����+H]�����˶���,/Pc��?@W��8�����b2�{������7��U�:�ƅf�H��������6�����+��w-���f*���׎o�|��Y�� �k��^��Xz�Ȗ��W�{N������~چ�sֱ"MT}���o�׎o�|��Y�� �k��^��Xz�(��¦�L\�kg�Ť����� E��5�O�U���.b!��u�w���v.���A�I�z�9w+�!J�0©	]�,�\DW.ɧ/H>y7�J�]f7\��1�T�g��������G2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcn��^��N�oߛN�N�FQx�0O>�Y�<]/2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hF^����i�̨���qh�'aba�	���
��?��n;�|-�Z��2S ���k��m���$[΁�a�n��Vk��w/&g�-ΘBdN�FQx�0O>�Y�<]/2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�tw:g�V|�hi��p�7��Z鎬�����R�LM��ħƿ�9c�1��8�h�� ����f�#�eM�f<�,=K�F~�?|�[_c9��*��OT��]S��f����om2�����iҢ��V�x��%�a��i�9�J��$b6�]ʆ�In��t@���z������)����")�^�3��8r�Wk�ǻow��R�nI�GI$��ǂcY�~遅��'�:��'n�^0o��S��S�Ib���ό���.ӥóM�˄NQ��臿5"c'��ɿ��3P�d�8!��vp�P}��O���w2T��b�T��xd�Y�I�;\h!E��c�G�*ZkS0��nB�+������]��)`���"��y�LN��K��g����R�<�W�C%c�����<�W�C%����_Wr��;���EWr�L{1��ox ������ �i7�sp>{=J���.��W�}�"�,�>E����\�vūx`��:��g�0�u�L{1��oxr�O΅��C?�D�s�R�"0��<��	��������JF!՟Ր��M�aW��Σ�?��<��z�"�~��S�
/P��Ѷ����A5wr�4�Vgn`��p���n�O�V�N�s
l���u���NX@��^��>��}� ���O%��y�䃶&f�����SVc�5ߧE4��?"����a�m���q�l;1�]�I�rT�8#�>-��;��S������yq]C
R��T
�N�oߛN�N�FQx�0O>�Y�<]/2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hF^����i�̨���qh�'aba�	���
��?��n;�|-�Z��2S ���k��m���$[΁�a�n��Vk��w/&g�-ΘBdN�FQx�0O>�Y�<]/2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�tw:g�V|�hi��p�7��Z鎬�����R�LM��ħƿ�9c�1��8�h�� ����f�#�eM�f<�,=K�F~�?|�[_c9��*��OT��]S��f����om2�n�h޶�\�Ji��'�o��Q$������aU��D�	a���(�E��!�`�(i3l0��F��j���^B_�(ba�7�X��)z�s�!�`�(i3%Ah�%4
>��XP��Ȱ�^�7^/�AJy���l�f�nϵ ���3�ҺIÙ=�H�}ʧ8Еb����������gE�,�Q�^�y�zL͊�q��_�0���ӨI��'���Z[A�E����F�'n�^0oL��pN�5����`K�x��R͖"�,�>E����\�vŻA�1�#`�͌4s+�ny���A�!3v!�`�(i3JHn��z� �&�^`(���%�a�N�+��#�!�`�(i3�b9���6,� k\\1�*_��hc�ʹ���`!�`�(i3l0��F��j���^B_�||�?�5���J��xi��͆'�X%Ah�%4
>��XP��ȵ�d��w����y{¦�$]\� ���3�ҺIÙ=�H�uoglR���c&;�p� ���S�Q�^�y�zL͊�q�� �-8���I��'�	�ų_��E����F�'n�^0o%|�J�0�5����`K��q��"�,�>E����\�v�Qq
˟6͌4s+�ny��9� W0�!�`�(i3JHn��z�k��%��6i��%�a�x�+Vv��2!�`�(i3�b9���
Ay�9�6>1�*_��h���Q��~��
c�[��ƣD��T�����NI�����m�2�Z,qC͌4s+�nycfl��6t�$X4P�JHn��z�S@�z�R3��%�a������?6�9������7s�9���o��S8��%�CF�I��r��Ȯ��ߊ��H�R�?�ɺdX�-�B�85���%�a������?6E�C�Έ��7s�9���o��S8��%�CF�I��r��Ȯ��ߊ��H�R�?�ɺdX��<�-���#�p������p:�2],˶�9�c	o'E!��s�Zu�EPD]�I���2�����Vc2�����Vc2�����Vc2�����Vc�
+&�s�A�F�7���3�GXS����E@��~���($�J.���
�=W�֯�^��N�&��?�2�1p���}������]�0�lK'���Xw��_
�u�m�\��q�Z˻r������U�r�}��}����ހmu�m����y^�k���%H�$N�oߛN�cL�qh�  `C�H��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!��D���X=��f��i��зq8�ЈxKʜ�#xI+r�� 0�D�A��t��D)��i�d��`m�¨3��%�$�������\O�a�|�6����&��DErwⳘ=�C. ��f?��s^�xct��_Tҥ!�V��NR0�����O�,�WNT�N D|�5N��VA}�v�a'����\�Z��'�Wa�L��ʻR0�˧���.�E����Fr<���\�g�-ΘBdcL�qh�  `C�H��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc.�
͹U��k�t���L53�����)-}�vPt�>xA�ꓩ�l;��!I/�������A��1��+�W��J�ݨg4$ _o����OI��@���:��F�b��@�zL͊�q��c�sYIJ8��OI��@�n���������Wq{�f��a��{oS�=wK��7�&d&(C�#�7#^�Vn�^ֻ����XP��Ȇ<�qp^S��j.Z��$�sӢ�]3�����c��(r$����G���'aOދK-\��$-��Ǡ٥L����e]�u�����!�M�T���ݏ��A�!�`�(i3���+�J�������"�,�>E��W��Ґ�YjZ�p��Z����r;��*!�`�(i3"�,�>E����\�v�!�`�(i3Sn<Z�)K|K�@�����!�+�!�`�(i3%Ah�%4
>��f���T,�;C@����%?!m�Az�F��O�4p���eq��VZ�0�s�b<�B�_���X�KM�����7������
�]qE�&���W����Q�^�y�����9�!�`�(i3���3�b���-the��戉Z�T!�`�(i37s�9���o��S8����J� �j��h@S�@�]_LO!�`�(i3JHn��z��x�f7﹏�1β��h����0���,�W�B�޹B$~s%��@�:�����xwƄ�{Ƨ\-TX�Rj�+s�!���r��*y�xDp��T�/i�M���"�,�>E����\�v�!�`�(i3y�Er�)=�ᏅN~z��9�{�G�K*V׹ږ��_��f���T,�;C@����P@zQX�76�$t8[��5��FX9�p�x^/8�D�n�ؒ1ECWI�R��R��=���b>���F9M؛��&�}�(�dW�,��(�a�肢�{l�f|�ό���.ӟ
�r��	G$��R�lD<��z��}�Q2�+�Yə~�yD݃��r��DB�����I�b}Ω:���V�(^��<��z��}�Q2�+�Y�7
�4�.�E����F�ҋX����|P�������A�=�8bH���L��B�;#5d���7Ê7�E�4'���Xw/���:;aR[�T�.�W���1�}�ױ��(@�E����F�ҋX����|P�������A�=�8bH���L��B��)�ޭ-�7Ê7�E�4'���Xw/���:;aR[�T�.�W���1��)$磨'jU-j�`�ҋX����|P�������A�=�8bH��Ę媌�+�<1(f}ظ{����$ <��HT� \r���㯄�����
L'���Xw��RN�-#�ьb2up,zk�g��[��v�$ƪ;���Q��/(A=�kX�*1�e38����2�9)�����m��T��J<�]qE�&�owђN�~R�wX�յ�8�,wO۳�yz�<��z��}�0z�cUL� ���Q�'e����u*w�A	'���k(�պ6<��z��}�0z�cUL� ���Q�'e����-��\4vߖ%��mz%���=a\�&'UR�q������3���R����o秾�!a�v�����w:ꮆ@IE�U��@�ڗe'a�v�����*� ���@IE�U��@�ڗe'����h+������E��@IE�U��@�ڗe'��;R����H���i�Ox�j�d�ƥ4�,�:�'t��t�W�lT[�HF x>H�|�Wǖg3ȓ8���/�A���0v7���V�x�O`�����
L'���Xw�j�7���rcJ]�0ݫ���Uh1�gؘC���t\>��fm��]2�y�Z鎬����)��e���Rf?����]2�y�Z鎬����)��e���= �J4��]2�y�Z鎬����L�`u�K�˱�Ui��Q�x��8�,wO��ٷ���TD��-�`��8�4�%��mz%���=a\�9�K�v`0���'=��"B��$I��w��,��xc�l��m
��5�(�����:x�V?W�)�ޭ-����
L'���Xw/���:;aR[�T�.�W���1���~������yf��?N/7G#+������z����A�b�*܋���ԓ�Dd�<�,E9|.���%�S��v���?�R����o秾�!rF)���X�3c/��!ő!XF3�@IE�U��@�ڗe'rF)���X�3c/��!�:GV��d@@IE�U��@�ڗe'rF)���X�3c/��!P;��	�@IE�U��@�ڗe'rF)���X�3c/��!4V(�x@IE�U��@�ڗe'rF)���X�3c/��!з���jf@IE�U��@�ڗe'rF)���X�3c/��!�f���l @IE�U��@�ڗe'rF)���X�3c/��!�Q��Y��@IE�U��@�ڗe'rF)���X�3c/��!��8�ۦ@IE�U��@�ڗe'rF)���X�3c/��!��A Ly�@IE�U��@�ڗe'rF)���X�3c/��!k�O�`c @IE�U��@�ڗe'rF)���X�3c/��!����4��8@IE�U��@�ڗe'rF)���X�3c/��!.�0�;l@IE�U��@�ڗe'rF)���X�3c/��!'��t#~t@IE�U��@�ڗe'rF)���X�3c/��!򊫖��@IE�U��@�ڗe'rF)���X�3c/��!��];p��@IE�U��@�ڗe'rF)���X�3c/��!���L���@IE�U��*�QN��� ]���f��v�鳔�Ċ��8���K(��z�j�;9�e��L53���Z<�~�q��]3�����c��(r�CRQ���E�+d�ίp��V�����Y����딼�\�v���T�©�#��l�َ2c�'z͌4s+�ny�X��{��ܛ�	�����^�%k IÙ=�Ho?Y���	3�Ð�9�X�e�B���<����ą~c�PƐt
����������\�v���T�©@���U@���:��F�����XuY*"�nw��F�dZ0o�v��CRQ���Eu<�.��	�L�t0{�A����8V�l0��F��j.��h��u>1�*_��h��Ӯw!)��&�t5C�,���m�b9������U.6����sd�Hc�.2��w�k#�J����͌4s+�ny\D}��^�y�����"�,�>E���]�!��	Ǹ�y85�|읯2�9�G�"�|��ߪ��wZ�n��[��rs�(�̴Y�{'%s�6F���y�8� �w� G�"�|� }�Ri.����l���r{����JDn ��aů�x� ���rs�i�H���N���w�Ve��t_-Z��T�\ ��QD� ��-a�vݝh�c�A�L'��KD����w�Ve�U�ԝ5�͌4s+�ny7\�%Lţ}���u=|�z�)�]�!��	Ǹ�y85�|읯2�9�G�"�|��ߪ��wZ�n��[��rs�(�̴Y�{'%s���A0�>�8� �w� G�"�|� }�Ri.����l���R�0�;"��9�{���|hY���rs�i�H���N���w�Ve��t_-Z��T�\ ��QD� ��-a�vݝh�c�A�L'��QV&�f�w�Ve�U�ԝ5�͌4s+�ny�y��P�p�V��O"�,�>E���]�!��	Ǹ�y85�|읯2�9�G�"�|��ߪ��wZ�n��[��{_8�Y���˂lq��r'��i�B�J@�l�s[�5����`K��D�	a���Ӯw!\�8䮨��ekW���I|JHn��z��ea���4p���eqd���w&�r��VYW\�����[!�`�(i3%Ah�%4
>��XP����~��84Z�Ћ�l�TE�խ������S�0ů�x� ���rs�i�Vw�C�-��0#�tC%Q,!�;��
r7��(*h�Qf�kCH`=Th=mP��T�͌4s+�ny\D}��^��ٙ�D�s^E��S�Z鎬�������(���E�̱!\Z>�
6������+$��g��U-�e�v�W�G�[�^�������-the ���mh.�]����GC.�|���~��H��efm�0z�cUL���a��<mDrW�B��"���PB[<b�P�`<����B��٥P5���rs�i�H���N��C�X<� ���B��8�R�Z_.΄x�g��	��S8��UV��\Ƴ�r��Gh�Qf�\l{�"7�sa�vݝh�c�A�L'�1�d��{�ʬ�缆�YW)��͌4s+�ny �Ǧ�_@f���_t��R��XP���x���: �&�(E�{�ʬ�缆P �8�-�US�����U[�[B��$�����˔b�7D�EI����I�O��\�v�d�jFB��]͌4s+�ny]"Jׅ����d��.%Ah�%4
>��XP��Ȱ�^�7^/��1������p�V��O"�,�>E����\�v�VNub��pzl��a�Ʀ�|þM��a��zr,/'���Xw�j�7��r��&D�:f��:F�X?�g��U-�e�^.�@���e��0�U+�qbp@���K�Q�f�;�>)ʁ���f��Y�{'%sgeߪ�{ ^�x~�(vi�t�c,�q�T�\ ��-3zYIިuIF��^~�$�x�Wt!�`�(i3���+�J��Y�{'%s���䒼�7��Hn#���T�\ �͘�f��p�b�z'hۉ)���	4ˣF�n�5��cz^8������зq8�Ј'���Xw��fi~�'K�2��J���"�!ɺy���B���Ȇb�L���g�"�,�>E���]�!��	Ǹ�y85����@�`�8�Wǖg3ȓ8���/���fi~�'K�2��JHm����v�V�Nt�s$]�6����ޤg��c�n�5��cĭ#�?UM�!�`�(i3зq8�Ј'���Xw�j�7����o_��ü~���U��g��U-�e��)���UM`���R.OƋ.]$�t_-Z��T�\ ����Hq���F x>H�|�j���Iq��w�Ve�!8���\/Üy�a
�:�,�!��qƸ "g��z�WCp}��~Ϙ�g����P"X����G�"�|����.N����=��Ʒ����V�3��yɶ7s�9���o��S8����iY��"w�z��C���g��U-�e��)���UM`���R.���b\�#@[�I��Bg����P�ߪ��w��m�C�7���s��R��һY~����j��n�t�q�ٲ��+�J��Y�{'%sAX���	q���b\�#�y�Ya�I��g��U-�e��)���UM`���R.���b\�#�y�Ya�I��g��U-�e%uX���4N�|��Z�<kx8냞�!�`�(i3��Q]� _Fr�����WF!a�ޅNA��6D���K�Q�o{��:��(�[�*��Q]� _�rs�i��O3JT�!I�T�\ �͘�f��p�b�z'hۉ)���	4ˣF\d�RI��������yبw�ሑa7s�9���o7�B�J���o{��:�N�#�@j��{�`��Ҝye��B�o�\q�߈q	���S�[N��t�$Z���>�ߜ�J����^�_�J*�(��Z鎬������D��찔q_�pk����2%g�#0~��}�� л��@(�Ϯ(����%��yBD~"[
W���VYLl*w�{	�C�9Jn�+��Q]� _Fr���������0�@�U_� ��*ߵB`���!�`�(i3�!��@y��=�-Ǻ�:Nɲ`wl�����`�Ǔ3zӲ݌���������j��-�n`5�fK�Q2�+�Y�E�!Up-i�Cߋp{T���[�2ٛ�X�/R��:2QYeƈ�c�Z�~E�!Up-i�jK�o[���[�2ٛ�X�/R��:2QYeƈ�c�Z�~5�e`��9d��l����v�}���X�/R��rs�i�H���N��/Üy�a
���"X��[�p C;8;kѶ���� ZkIb!8!�`�(i3�d�٣�����6>�����ev.������f��gy:h+i
Z鎬����Ĺ#{��a'�<� \�Q�w���*��_?�v���Q]� _�:2QYeƈ�c�Z�~ݓ��E�I�Q�Тd�!�`�(i3�d�٣���,�JL���+ޡ)Ծ�/�n�*���?�#�6�fȯ�?
YT'���Xw�����C��'��/��࠮R:������V�6IWJE�r���秹��ч����=ў@'���Xwd�n]N�^ �7�}3��|�b�@a(􆿳���Qs��������=�8;�(�[�*!�`�(i3Ww�[h�q��!���\���Ȑ�'t��t�W�؏ 4�+�{_8�Y��M��)=໺(ӈ���x|}�|0�(�Y�MM��5��g�g�(�[�**�k�����\F�^�	E��߅�'e���婣	���U�dN�<@Iv�H�_��Q��b�z'hۉ)��!��|"/3�+��m\ƪ;���Q�0�=s�����[q�2�ߣ/s����.Y�[&���,�v����z��ˇ�h��ܙ�[-<�+�my$�N��YͲ�pzl��a��Ǯr!�`�(i3!�`�(i3�n`5�fK�Q2�+�Y��׎o�|���Y����!�`�(i3!�`�(i3�d�٣�����6>��i�X��*Z�!�`�(i3!�`�(i3�E����FZ鎬����Y�V��#qFL}��!�`�(i3!�`�(i3���+�J���q���U�pzl��a���gE��҂ϱ��[��Q�#<4^��n`5�fK�Q2�+�Y�kѶ���� k���3�F�-XX!i!�`�(i3�d�٣�����6>����9וP�;xB�_/�1!u7}:�E����FZ鎬����Y�V��#q胬<ċIX3�A���\�J2)V���+�J���q���U�pzl��a���gE��ҩ���;//M7$����n`5�fK�Q2�+�Y�kѶ���� k���3o=�<*��e���b��d�٣�����6>����9וP�;xB�_/]k�WM��q�E����FZ鎬����Y�V��#q�?�B��{k���3�z�Q�q���+�J���q���U�pzl��a�-{�*�;�Eo��K��]�q��n`5�fK�Q2�+�Y��׎o�|�8����|�M��5�!�`�(i3�d�٣�����6>��P��r��c� v?b���7;�Eo��K.�wK��� Z鎬����Y�V��#q{��>]#���)y(�O|�M��5����+�J���q���U�pzl��a�����;kn�P��l|�M��5��n`5�fK�Q2�+�Y�K=J��(��I(ީ���a41h���������d�٣���Ni�4�ڼ�t%>^��?�y��hL5ӥ����c^����
<ڑN���2�A��1��R�9*�eaA�|j?�d���&���>E��*�(��z�¿-ǂ,yߊ��b,�a������)�}�����T��.��W����t�.�!�8�}�\���;A<�SNp>�3������"h���ƅ5����5�`��N�W'�o����f7����e��x����#E`D���$G�	P��?[@S�CZ�~۵�q�#�p�	;�0�e�n�xdɨu �䆡X�dr�jf'��H������V���
���F:_ʣX`��_/��IC:GMG�2�3�A�E'����>E��*	Z�~(jm�7jl�N�Ar�/=�N�}���X	j�w~jiǎ[��S��_�:�R��h�4�b"����gE���Y(��	Q��H/!�Sy�+�z�}�-�%Q�a�4f�+�Z�{�b7�-�4T����	��,��<����r�k�,��~��U?'�����ٴ��{�G��ͫ������:[ۚܖ��`�[�	2�GF�&���#VW�GaAO'��7wT�,���P�&`bH$��>��L��$�I��i�j~>�Q.Ss�@�������-R�X��%�VB�=����R��(7�
��o��N⃟g��|"u8��d�w(�`��l4���/A� e8�~��f��Ԡ8�tF���)e���n�`�v�Q��7[32X|��h�ɑuϢ\�S&��)Q�����{1���	m���N����B�c���7zxs�ްs���	m���N����B�!2^D�S	�o�7s�����-���
0yS_,D]8@U���H#��Ɵ���X`.�	����Y�oc!���ٴ��{�G��ͫ������:[ۚܖ��`�fJ�WM�.�A<�SNp>����AnJ��ó)�󼅯|��%6�Y�JDFH��z���8�ϑ��[���D���0�j�J�Ñ=��[1�%n�@��V�����Y����딼�\�vūx`��:�,�qo�,ܛ�	�����^�%k IÙ=�H�]ƭ��&d&(C�#�7#^�Vn�b9���sW��NZ�uw�@.�/wc1��˪Xk"�,�>E��<��z��}�Q2�+�Y��1S�����Y%T��BPS�)37J*u)T{6T'�f�;�>)��U֔�>V	�]�!��	Ǹ�y85�R�m�.wa�Iz#1�<Td��"X��[�A��N��|�+�� VU+I�z�c�5����ݱ�Ʀ�f�������~T�����A���gf׿���$	n��s��ͫ��;���^hq��:0k�y��HzL͊�q���19TH���8�6:�F!�`�(i3l0��F��j�
����uK9��>�������q�}5h�-tQ���͖n!�`�(i3�b9����6�{@$��uw�@.�/wc1$�W��9��I3���S�)37J*uc�A�L'�	�Vh�/�owђN�~R�wX��v~S*��R������5	��]�!���������RP=	P��{l�f|�ό���.�L�2�r�Ĳo  ��]�!��V�,�q^���ȍ�)0f���{l�f|�ό���.�V�|M�������5	��]�!���sC�)�.;�<.��{l�f|�ό���.���S��"B��$I��w��,���|HH9M\��e���S������
�:�e�ӎ�4���S������	�_���X���n�k�r�>?le��pp��]�!����-joG�j��ԁÆ�7G#+�ǟ
��|�6�E�W#��e�0
A����l_�U�x��3����Hhqu!���5�Nn���4L"�#W��xW�Kg!�h�����7�$�G�j/����X�e��}c���G��m\Ӓ�qܛ�	����(:��=�M��0�d�Sd��_�a���n�|Wg�|bVzN7	+`�9
EMܓ���;�e >���l�n�Zl��Ͳ�8�3
�{�-�>��t��ԱͽP�nT��Э��y�L*���8�^�.eO��q��S��;�(e)��v��=����'�$��u,��y�"���Չ-d��r�b+��/6!��Ei�gz�����n�|W;"V7��evwJ���&�o�\,9o$aϛ`!�A���
+,I�2Sj�	�$ɜ�\�۟�-?�d���&����{ԕ�h7�{`��������* -��ed.:E������ƄH����[��2����s�ZK5U�㶰wi�G�A����`�+N'����)�!9x�����A��Y纽|ԯ/��m�h@ѐ�ER�)��<|+!N�e[�������C1�у�ӌ���qfb�B�l�2�����^t+����2�\��v�"f$^���\�}�J2)V	^�����v���?���1S���������;q&1f9m�҃kG���!l!�`�(i3W��N���;�������<�K�kσ�a��R�#����[��G��mO.�����R����ć��mRiP���uVw�������`�-<�B<.A���0v7��)�ޭ-�΃$%HJ�#��|�k�HB���15�-�bFd%��I(ީ������	��+?�d���&�Ա��+��i���%Ὠ���0��H22��=�z#����2av����pJ�B�	e�q'�D؉��_�m�����W���9�b�w�䩳J �s���H@�{���]K�I[;;v�W>�.�5�O�O��S�7����eߖG
�<ݬ�K������,����k�*�.�a�n'�,+$\�M����F�V����Z����H�ЫY3EZp��Ĺ� ��p[�ٕ����se�{�z��x� ]
�"ǩ>�)E���Z��v~S*��R�J�a$�Y 	�z��V��2�jE?d�1S���������;q�Y�f�ƥ�d��Ke�ά@�ș�I����~u�B�f��.X���ֻ�����h+��
!O:0��O�W�."��ђo�N����C����N���&U2�S#:�*a��E��]n���G�87�]���`�-<�B<.��U4�i%���;$�{�R�$�V�o=�<*���Nm�}��0����8�D���"��	���Yb�V��	��y ��f"�$�!����L�����©h\���k�9�����/	è��0�	+�����6(���j��h@S�@�]_LO�Ŵ#����#g�k��m�z5�Ւ���Z	L�'�}5� }�	��%���K5U�㶰wh�(R;�����3Y쐅�	|�Gy0E��*����	��۽IM>�������ܪ/���ܸ���$�;�5�sw���J2���;B����ՑK�^��F
f����w	}��tsb�?r	�'3���EK�����
�F���LS�ߛ7�C|�L����5uE�(��*O)�J�1U"��2 9�Q1~����?ON���?�� 5傟������kV�U~�X��9&���=/
��G�~7��|YYp��]��nq/����[΂8�:b|�%���,���D��\��%��	��<�T?N�·�����9ۇ%p� ���3�y��9�<�{Pkt����^�r��3�h�|��4-�Q@_8X��Z1~�g]���f������y	��Bo���+�hi��;	�v�鳔���bL�%s�^�� �	���bl�����7�-m��0����NF>4P��)���=E~���e����
��M+)U�D���ڡ�$��2H��&Y��V�'��С������$}%��oR��ן�/��-ށ� ��*lxi#�3��|��4-�Q�p����i�7-ڍ�mI�ｘA ��
�A�m�`�H_�U������%Ik�cIƼ̰�m���;��u�(�};�1F�]�q:�q���8̈�f�������,�Ȍ���\�H�f"��ɔ!:����kݛ�l�a�t]p��Ү��~�[_.H P��?xA4����2��<E눏����ܪ/���ܸ���$��L��ߨ����f��C�쌓���2�����=S�vʐ̡�&Y��V��� ���)���F��=��'?$���0#��=�\���@���,2���!*�؍�~X��a@=�����Yx��t*�=a{��67�M��(�K!2�7�&���=R��
G=�H�쭽�o����rN�>���t�'%��H��܌z)-t"wdC��_m+ �����*��W�Kb���Z��KD�И|��,2|�Z�F_u�
!O:0���.�Ҭ�^}�]���k���3�F�-XX!i�N���&U2������PG/�W���LU�L���)�lV7�]���6��(�N�3���?�xB�_/1d�H�Zc�{�R�$�Vִ��l�+,@�uU� ��}n�8��D,�K�-)K�'h��Q�C��1Dm@<�9�X3�A���\|u��W�s ��9�Q�Z^ >�@�uU� ��}n�8��D,�o�fy'h���I(ީ���x�tO7����[�����|\���sIN�vvH����k����ɝ\�!2A8�r<����P ��BP�wb�H�Z�^6w��<��D0m�'1{{!LU�L���n�Zm����)0kcj1�kD�t�Sj̆���K�|�'�ȵ�]u(+֢���S,�D�c��Qԟ��
�A��R�j`D�����4m���Wӭ�6@ri��P-{�*�;�Eo��K�p��h׬V�!+���}9��m;�n�i?3�(��'t!���Ci嶨��V����m�=�er߮�Ȗ�%T#�5��gE�����b�ђا�0�)_��c%����lxb�뤆�J�e�C��1(�����d^_�Rꑽ,�I�d�N�1�b�*�4MM��Hi嶨��V����m�=�er߮�Ȗ�%T#�5��gE��Ҁ�M����]��Y;�c%����n������И|��,(�= \	\�M<̜Z���wt��B�A�M�I7g����i嶨��V����m�=�er߮�Ȗ�%T#�5��gE��ҩ���;//��0�)_��c%����yg��c|q!И|��,(�= \	\�/��������Ch@�����y-�c��d��ȵ�]u(+֢���S,�D�c��Qԟ��
�A��R�j`D��R'�u)]�t<���J�?�� w��l�iu��T�U9��
�;�Eo��K�p��h׬V�!+���}9��m;�n��(��H��_�0��R���־�U��sp֟kh�W�f����C;��҇И|��,��N�i��!��z�w��<��D0��8#���#����a�9�;�Eo��K�p��h׬V�Sy����!�`�(i3w?�W�S[И|��,"��7Ch�m�1S���������;q-{�*�;�Eo��K�g&�?�U.;�<.�����^��1uv��e���%�G鉖�;�j[����"��8�O_���`���k���3�˙	e
^�I�*�y����(@CPwn������И|��,"��7Ch�mRiP���uVw�������`�-<�B<.�,�I��
���Ƀ@tl��(Ur|u��W�s�ַ
���iW�\G���J�e�C��Lle�J��0����1�T1���T^���И|��,;�L�����G�Ȧj�v���� έ��F��#�Ц�w�L�������"�$�㔩?'�m�6X���(��ޭo:��gڳM뵨�I6�j4̗��W;��"r뾃	��s�Gq��M�B���޹B$~s`�� �:Ft�EO�{����O�2��a��x))b�K���$73���'���)E������?�d���&��n=:�Ed~z,�	��lx��`�+N�%'ף'���i�7�^��X��=����`�+N'����)�!9x�����c6�c��A>	�x��FR��GN@����x�hn�B�l�2�����^t+������\��vMjm�f����qfb�B�l�2�R"8�{����=���z���X�v�J���C�O��S�7���޴:�Q�� +@����T���!�
���qfb�B�l�2��e)g��nQ�4V|M����io7�N����qfb�B�l�2�R"8�{����=���f�H�Γ�^���\�}&�1d��̺Eh�m-6�c�����0�J����<���r�G���6���U6!w����}q����߄1�9F[0�#����X��=����`�+N5|hy	$��EV_�[(����R�?d������?���+y��"nF^�{��s^��I�$nx떖ݏ��A�7���?�!���bJ���WW�+���3��0��A����}�ʩ�Vh�l�G!W�:4'.�Rי��3��0��A����}������T{�o�����'N U����k�*�.�a�n'�TJ��H�*�b�>�F0rv�J���C�O��S�7�����)z����=���f�H�Γ�^���\�}&�1d��**����r|�>��B��;��|B������CU�G���6���U6!w����}q�����_[�xT�oH:�m>@{'���da�v���ޚ�^l��{b���g�1>���A�� �8 �\ �Z�����Xe�����"��]G�PG{��_����0���p]DWl$�`�]
���blm~H�+,����2�����~y7�`�9�O����۞h�G����M�趧�,�qm�c�,�[`�?�{�2����;�H���o���6G4�?�C<xWY�K��e�Igg�QuU�����DZܤ�j2t�ch����	'����'�SS������{�T�`NR���c�,�[`���O�:�2rF)���X�3c/��!p�=n�٠��f�;�>)�L��<z2���	�i��#�f�;�>)�|(�כ��	캧xӍ.�*�yȩ�,�+KK� ^���PG{��_�����*�U	=Q+����]
���b�/�4e�{rF)���X�3c/��!�&�?3o_��f�;�>)����k[�R�<lͬ۞h�G������W����I�&�`���Oam�87/	��ee�PG{��_���/�>Y�]DWl$�`�]
���b��R��3���2��h"r���Ez	*HD{۞h�G�CŦ�KT����,�qm�c�,�[`�j�a\�����;�H���oCO2��?'?�C<xWY�K��e�IggI]eLu��DZܤ�j��"z��U��L�(�rY��'�SS��yӕBn���'n��c�,�[`����R��߶��,�qm�c�,�[`�t�U'#�;�H���o�����jw
�q8*�n�5lY��fZsdDH���Z鎬�����LE^��EjsdDH���Z鎬�������(���	����Dj�d���m����0+C�t���� ��/��}���.��s��,��+U�HJ�h>A:����������O�1��`�^Y�{'%sAX���	qOƋ.]$�t_-Z��T�\ �̈́��L�)@R\�N���a6gBa�����0�]�!��	Ǹ�y85�΍y� I�M{[���G����"X��[w�o�4�n3���+}��l�&�Yw_�����\e`,9�H�W2%�ܚ�!��@�YZ[4%|S$N\l�IQ2�������C 1]qE�&�.}�I�̆�U�J�J�ƪ;���Q����Cs�O� ��:y�;�7�E���{$?��z�(�V�ܼ��Yu�mVNjƪ;���Q�+ج ���k������������9��*(!�~���i�x*vX¸`��;R���\`o��ӎ<i�LE� R8�k��z-�%��u��;�j[���.��o�܁#�s���	�!��n����[�(���u�F8O*�E3* �s*F x>H�|Ċ9DX��&{H�3)-(�K��*���@Ph�9�(P��a6gB9��xQ)?�NjX�U��E`����(�V�ܼ�ʽ��φ��<�6��ך�$@-w���"�uA}�/��4�磕�9B`�n]
���b�L0J���g�0�u��j��W�&�+K���n��A�ԩ�x{^4��*m�K�"A���.���G?�dN�<@Iv��nt=:�6���OB\����^a����HŹn�軑��r��4M̍����;�H���o4Go�HHm��1��X��WG �� ���K%����	x=:���	�ج��	~p�ܩv�~�E��z�WC��"X��[y߉�m�$x(�i��/Rh�x#�L_�(D{ͬ�y�4����gSS�[nl��#� �%"%vv�J�ԜM����}{}�z�����v�Y΃xI��o��#o~��H&���'��N��i��x�l��15�r*Iީ��>��yܛ�	���n������7a	����"���P1�߽K}��[T�)������x��\P�O����X�e���&qL�+.�/'��Y�
�n�5�F�^hq��:f��3\z�[
�}3��*���1���v~S*��R�-����,�Ӏ(��c���9�L(�y�}�b��H���۞h�G�֑�t�ʂ5z�¶2������텙�Cߋp{T��c���,�\��{ElCg?	��ofob0�۞h�G���w��z�=k�Rm���8Ơ4�ܩ"۞h�G���7?7��R*E���&�j!�\B>�jK�o[���[�2ټ�mˊ��ձΐ9xWW)��~?R����I�
�2���L����\9�oA�d��JXl'�&�P�2�PUг�|<�ɐ�>8�co�v[�(!쥭*����	D~��n�&�;|>r:w�:��er?G��7Wx� Pabݙ��N�g�c�`�ɐ�>8�c�"�rZ��.�uO|&�9�r�I�;3�p
��a.��,	�g��WN������)<�-w�|��qĵ=)�7��B6Ji����|���!9�j�m�����N��4M̍����5Ɇܾ�]��	He)O,�rە�f�;�>)�-m>c.��{t�Z��P��3�Q#� :a�	�+4D@��/�ciJ���z 7	B>�b��O����~y�
3��0�ǳ�ȕ<dh�}3d�jK�o[���[�2�֚���,��Hp9��Ԍ��Ǐ�c���w�I�7ݟ=�NM���ɛ�?ө�&�(5�;2�@�a�����be�vҜ��)P�N�g�c�`DE8k �Υ4^��)�d+�����q9+t�}f��1�x���~?R����I�
�2��f��U/��.�[ ٓ��r_��mԌ��Ǐ�c����3�6oݟ=�NM���ɛ�?ө����h`�CgD�|�݄����Mv!���xx(�i��/RŻ�&ǥ��a���F�LFC7�5$�)�vx/�k
�SR��Y0R�ne�>�H�ܕ6��HHD�u���&.)+�ޅn���(��h�*蓱Wxi��o�bB�۹�D����=��Y��RJWz���
9�5ARL��׿"aj$�b�w}P�
���(�����d��R�Q��=�ƆR�(o�Y�f���'v�qB���jK�o[���[�2�gu�}���<�f�;�>)�-��a�A�so��%���;�N�cP��&��h����E�F6���Wz�o�3p�60���!��2��J�J����3%E��_��=��}xsEqFM���K����x�l��15�r*Iީ� �����Y~��`�J��xG�"Dd&(C�#�7#^�Vng�m>�`^����S,���� w̭T�&��is���'��� S=?l�_)��~�b������7ZON.N�N��;�Ż=qW�e6!�;�H���ow3Ԁ;M>���4����τ��;�H���oU�4{��F	��`i�8p�u�$��-vy�R�QY`�CgD�|�fSr�P�
ح+��&�.6�L
̸#@#$Kb�i�bn�Ź]{?�����f"��0�(\P"F0�4�fՁ~>���37��f�������!9�W�Y�i�� �U�z����!Qr�g?	��o`
��3�l�g�0�u���^a����HŹn�軑��r��f��}BɊЇFH�N�u�)ֺ[�`^���gmz8>���_���׍)@�\�����f�;�>)��*� ���͚wS.6�zB��݋�^aw��Xái��ċ�!-M�O��~�~l>�.֚���,�%][��"��4r��)�N z�@�^�c�Z�~J�1���۪	�}a�]�w%�oφ��<�6�;�r1΀��t�e��99kU�#����	�i��#����UN�M��W38�G��4�V"s�ֵ�_%Dό��סزN� �w���zF������?M>��^J��3��a���Cوj�~�4v!4���X�#A�H��~?R����I�
�2�=�@)��۞h�G�jryX2�uso��%����,����«?�z�3$Ȋ���yu�R*E���&�Ut�\�I5Iy=���A�
�����ΥT�tT۳�͕���ָkd�vu+�vW�
�%��v��rw�&�z<a��N� ��M�W8߸��S�Ȍ��p|�
M
�q_�pk��A� FpA}�/6�o8:4�Ԍ��Ǐ�c���w�I�7�V@BɇF����������.gZP=�����p�>�q�M�4�(��o/��lk���t_��� v���il��l�=�����g-�B'Ő_�)!c���~?R����I�
�2��K�f�-M�O��~�W�{OEׁ��U_� ��*�Z����jf;[�������g�Z��3��a���Cوj�~�4v!4�����2?��.??�#�6�f��.���-M�O��~�Ѩ�f?�R���%\��o.��p*����H��efm�0z�cUL���ޤ�Y5x���:����S�>��a-6�Da�,2�C���l�yi��L.bC����f7� �/4�C�Ȧ؍�a-6�Da��0l���SZ��T��B--��cKE#�}N�3%�}�Kf��"������0�e�Z��j@�4Z��՟��G�0��[k�J`�\A#�ͫa���I˒��M���B�:����}7�������\�2���.Z��'���:��KY�[b%Ɨ�W�{OEׁ��U_� ��*�Z����jf;[���rw�&�z<a�4�ڈt�[b%Ɨ��q�;���a*`�(o�l�V(�ςMv!���xx(�i��/RŻ�&ǥ��a���F�LFC7�5$�)�vx\n�ޱ��H#�ͫa��R9�����K����0+C}f��hq+��=k�Rm���<��=���jl�iYX��R*E���&��P�>�n5j�?�T�^'��s_ㆂ`Z"�A(sB.��Hf;[����q�;������\�2���.Z��'!�`�(i3%��v���\�G�����dc�@z�ׅ�ؘ�X��WG ��\�,h������v�}������Ja�vݝh�c�A�L'0i���crp/Üy�a
��ү�+ҋ��/�ciJ��"|s8`69���TLB������K��"h�]
���b�v���V�i�;�H���o�4�= w
��ݔ��������@/��r �a�<d��]��9��6�j��n	Y'F�0!�P.	ƒ�3^�ԭ���d�n5j�?�T�^'��s_ㆂ`Z"�A(sB.��Hf;[���Ĕ�.p�1��zB��݋����f��)�F��2p "BC�I�#�ͫa���n�e�[7�w�sB�ƓX�H]��9��6�j��n	Y'F�05����Ǐ�{�`��Ҝ\ �k4N�n
V~$7���.L��h�T�D�ԗ�CW	�h9<���F#P�j2E�?�o{��:���m4��0���f��J�a$�Y ��\bʏq�2��Kk:)���2�z�X
3kZ��&�(5�;2x���'RFt�T��,���}��֏i�6rT�Xk:)���2��N�g�c�`k�J`�\A#�ͫa��l�Y��QZ���$#z�*�
��Gk>��Mv!���x7���.L��h�T�JDn ��aP�d���� ��U�_:���:��KY�2Y��+rB�0j�䴑f��6�k�*x$6�	�@�Vw�PV�q�-n
V~$7���.L��h�T�D�ԗ�CW	�h �ҋ�;#P�j2E�?�o{��:���m4��0���f��J�a$�Y �c�Z�~�X�H]��9��6�j��n	Y'F�0<gX����"�0S�l�%�z�J���o{��:�N�#�@j��{�`��ҜcZ�����c�Z�~�c*o��ܔq_�pk����2%g����<-����R��n5j�?�T�LW�_��%3�o�:�>je`��@d:�����{~�o{��:�N�#�@j��{�`��ҜcZ�����c�Z�~�c*o��ܔq_�pk����2%g����<-��ic)�̩��ɛ�?өx(�i��/R#k�˟ܒ�o|k�Lb��˓#���@�\����Ԍ��Ǐ�c���w�I�7<�	+�	�u@���kJ���af�iβ�=&��]
���b���M��#l/����1��X��WG ���ɐ�>8�co�v[�(!�,|7�_J�Ǉ��k��ߦc|n������$���h�T�D�ԗ�CW	�h�d���^�q_�pk��=��hX��9�{�b�o��/W�{OEׁ��z\�Q��TXP�e�g�6�<+s�q9+t�}��Ǻ6�(c#�ͫa���n�e�[7
$B�>���I����~u�o{��:���m4��0�g�F}kQ1�#k�˟ܒ�o|k�Lb�5ߧE4��J�1���k_���b_!2�͞nOY��/�eDɄ~����p���=/�`�&�;Z�MXH���3���~*�o��G,8}�;?�~�0��{�Zx���h�E�U<:�r�?��� N��r*�S	��5g=�,^sf�f�+�9-�i"'���Xw�j�7���sB$��#~��U���Yb�#<��7�}ퟐ#Â��&?�g:ξU64%��v��J�1���k_���b_!2�͞nOY�Ƹ.��v�!�`�(i3 �=Ú.��/�3Ĥ�!�`�(i3_j��u��[���MooM!�`�(i3�K���I9��A]ïi!�`�(i3M �̦�P�c��f�.E!�`�(i3!�`�(i3ZSX�esȸ�"rR!�`�(i3����ȇ��l*�����l*�����l*�����l*�����l*�����(��p�Hkq5��;��wD�w?⨻!�`�(i3����l��kx8냞�!�`�(i3!�`�(i3��a77�@���]�U��!�`�(i3	Xv��#E�l*�����l*�����l*�����l*�����l*��������~q,�!�`�(i3Q@w�ӏ{!�`�(i3�n3z(!�`�(i3!�`�(i3!�`�(i3���i�>�{��]�U��!�`�(i3G��0<]22�����Vc�R�
D~��2�����Vc2�����Vc2�����Vc��ɖ�~k�!�`�(i3Q@w�ӏ{��%\��o���|�[1qR���g���ȃ�ZK��������i�>�{��]�U��!�`�(i3G��0<]22�����Vc�R�
D~��2�����Vc2�����Vc2�����Vc��ɖ�~k�!�`�(i3!�`�(i3���dH�L��(���n����y��]qE�&T��Z=���i�>�{��]�U��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3T�����?!�`�(i3!�`�(i3!�`�(i3}S���2�����Vc��U[+��2�����Vc��f��w��]�U��!�`�(i3!�`�(i3!�`�(i3�)V��s��]T+�krB�0j�䴑f��6��ȹ�!�`�(i3!�`�(i3!�`�(i3��I�����6�|�MX9�G�tk!�`�(i3���i�>�{��]�U��!�`�(i3!�`�(i3!�`�(i3�R�
D~��.���{	RK2�����Vc2�����Vc��ɖ�~k�!�`�(i3!�`�(i3!�`�(i3��n��`
H/Üy�a
蟸���th�_ME�v~Aj�}-i #�sq�G]�K�Sb6�A�e�r���b8#۪��������`Z"�Au,���Ex��N�9�?_��s�֙��N�,�; e�=�#�vG"J�CJ+T �o��_�R�wَVݳA*{�;h/�0h�5eש�y�k�A�$����@/��r � L�#��e�wDJ��dN�<@Iv��nt=:�-���)0�ʂ�j�Ï��	�Li4"�	��z��R��Y"�g�YZ6��HHD�u"�T�B�Z�R*E���&�Ut�\�ً���N�c�,�[`���W�XN=7�}|��	��a-6�Da�����a�#�ͫa��l�Y��QZ���$#z�*[T�k�r٪@/��r ��%�z�J��\�,h���]�Ϲ���6�|�MX���%-4ɚrs�(�̴Y�{'%s�6F���y�q� ���+�6e���mn
V~$�u��XC��5Ek>2맫�?��_K��ⅴo=�IH�cT֓O΄x�g��	��S8�>���r8j�g����P�A��i������Ʒ����V�3��yɶ��9�W�"7�cL���	Ǹ�y85�΍y� I�Mkm�m#�m�e5ngY�-M�O��~ӶC$�-��xM��R,�g�zSB�������h��}�mT~1�����(��(��?��_K��ⅴo=�I�������3t���=�4�04�jf���pP�h�Qf��,2�C�����d����vk�iv��a�vݝh�c�A�L'0i���crp/Üy�a
��ү�+ҋh�Qf�}���ED����%\��oQ��u��e��H��efm�0z�cUL���ޤ�Y5x���:��7^���]�vv��I�����j�1>�+�9-�i"'���Xw�j�7��#�@(14~�����-��t���n
V~$����$[�ĭ#�?UM�C���a[S�.�go��8�K����ꪫ^�|U߳\�������n<+�1#P�j2E�?x(�i��/R�xȀ��D׏�����M����$[�z^8��)P�T1=�#P�j2E�?n����n���/N�b-�LLJ�|�HA�R��뛶��I��o6x�����&�(5�;2�f�;�>)�ӔuP��N([��}qn
V~$�A�3)]t����W����L��H�)l��T@��~�`�����e4^{�_��1��a"�!K�2��JHm����vx�*aE�P�HS|�4�04�jfJ�1����ݾ-/�uu��ڿ$�)�vxe�zA��;��|B�a��c��i)��]��ⅴo=�I��=-�!�^G�*$\��j��ͽ&�^������y�&D�H�B����1kܲ��b��\s��9�{�G�K*V׹����R?�d���&�t�d����6=J��}�7D�EIdQ�;{�r6]����e�kCF�(��4p���eq�x��ق$�E�Ν��J���(_\�^?'qKy���\N}zp�jN��;6ˆ4���Mt.K8��T�{��ed�s����y���uLK���������C�i�'6c�f��kq4s�a���d������^����g9�h�^+������������9�xV��	~�`��������!Qr��zj7i�j�}f��hq+��B� ��~���4M̍���kU�#�����1��X��WG ����Qj;b�J�3���y�my$�N���Uە���\�G�����dc�@z�ׅ�ؘ�X��WG ������F��Cߋp{T���[�2�|�P� &G�N�g�c�`�9�d�L�:��er?G�Wq�`ASi��ċ�!-M�O��~�����$[�ĭ#�?UM�C���a[S�.�go��8�&����vE7�MWO�6�c��$1ݮ�I�C��,�jK�3��u�!x�R���- ����%7e6����k�'�d0�(_� gg-	�\�G���:��er?G��g��ǻ�Ji��ċ�!-M�O��~ӿzR���b	;��Ǧ�<z!N]����Y�1Uj�|ᓆ�~_Nv���å;���.[r�gc�JV����l P�7��Hn#������Uh1�z�X
3kZ��5ߧE4��p�-a�D͢fU�9�׏�����MFi��|ր���5V��	��yx�_uE9�{�����ӵZ#=D;r�R��x�K粞ƿ��A�qL2�cR9�����K����0+Cd��y5\ N��r*��L�4��j�Ï��	�Li4"�	a�Xi��:��er?G��g��ǻ�Ji��ċ�!-M�O��~�Vb�ͼޘ&�jW� �=z��k�8�W��]���s�� ������uS ������)Ҩ�X,��'�J�y��˓#���H��$�W<�&�jW� ����L���ݾ-/�uu��ڿ׏�����M��ܐ�}�9Wi��p_#�����!�H��3�L��b8#۪%r�^0VEF�ߏ��8&�|��³ʂf>x�:	LtN8�,���	�E��zj7i�j�}f��hq+��B� ��~���4M̍���kU�#�����1��X��WG ��7O��4'��7�OT�,�rcJ]�0�{H�3)-��g��ET��w�/�K7͍��|��W&":D3
ڱ�Nq��5��g�g�$*T`�̂�nF���<�W�.�P��c3�fF�5.]����s��U;4���^a����HŹn�軑��r���/�ciJ�Kr���щ���ӮvZ��S)�3=7�}|��	��a-6�Da����b]
���b�-N�d�@/��r ��%�z�J��Kh*w��=\�1y*ط��w�44C ���8��9�.�`�ז����p�^ ���}M�ջ�3Z�(��{�vE7�MW�+�!�صzB��݋����f��ʣ��M��x{^4��*m�C$�-��������!�Lz��q�z=���R�����M�<*LF���i,��fx�W��L�rw�&�z<a��r����&�(5�;2����>q��A
��z(�����N��۞h�G���=�,Н��j���J�������ۧN�g�c�`��L�ΪA���Ǹ��St��h�T�JDn ��aDQ��;�x-M�O��~���L�ΪA�%�C�5��#���+�9-�i"'���Xw�j�7��FZ����^��h���LX��WG ������m���7�!`����=<�HIl:)�xq��44C ���(w"<��J!݉�����M�������ưCv�JDn ��aeGfFXջ�}E}��3��L�ΪA�%�C�5�ɇ����>�b��O���ưCv�JDn ��aڲc�`\%h�Qf���g��E�@*}��͖|���yG~Fx�W��L�;�#RՔ���5��g�g�݄���(w"<��J�=}Bnw�I e8�~���5ߧE4��tTi����[b%Ɨ��l"�$1ݮ�I�=}Bnw�I e8�~��b���e��!��4DE'z:�m7F���D�d�	y*ط��wZ3�z:��ˮ�N��rq��Ϙ��	�@�Vw��`��ZJdZ0o�v��%�z�J��R�����M�<*LF�o�HT蔊�cٰ�Ž��v�}����6S ��x���'RFtx�W��L�p�-a�D͢q��`�LW�]:vx��3AE�p|�/�GT�)�[�=�({���*Ȣ?u�J)':�L�p�^ ���}M�ջ�3Z�(��{��xȀ��D�[b%Ɨ�Ѩ�f?�R���%\��o�z��G�S٥P5���rs�i�Ǘ$� ��������-/J�����Ut�\��l"������3Y����Q����ۉy�T�����j�ew�]����z�,�X2���tTi���׏�����M;�#RՔ���5��g�g�݄���(w"<��J�=}Bnw�I3t���=�4�04�jfrw�&�z<a�4�ڈt׏�����MJ�1���۪	�}a4����@[�_zβr��S~��#�����!�H��3�L�N ��HdX�Q�����X���m����� :�>F�������f��ނׁ�4^����R?�d���&�(�h��E�3$���K��6�o8:4�;8I ��*�n89j��<$�g�0�uM`B�Ӑ�>�b��O�=7�}|��	}s�-���`,9�H�W2%�ܚ�!��@�YZ[4%��P�P-���F�Hj��b_X�XV�b�z'hۉ)��R��삍(�V�ܼ������A �k+Q�h'�Ȝxڣ9�$����3�� �fWT
Y��%r9���TLB������([��}qn
V~$2�t�N��Y���@�}%@�`�4��h�3��'c�,�[`�t�)
W�k��
�!���i��ċ�!-M�O��~ӿzR���b��C����z:�m7F.qi��rW
��t�B1�-�ErtI�2��i��"u���Ȇb�L��B bb���H��efm�0z�cUL���ޤ�Y5x���:����S�>��a-6�Da��g��E�U�!����R�c�Q��Ȇb�L6<�C�-�q���=� �������p�-a�D͢q��`�Lx(�i��/R#k�˟ܒ�o|k�Lb�5ߧE4��\�ܢ��,	սL��$����,�ǰ ����sԣz^08�2�# ��jߪ��b��@�)�H"�L��p�>�q�M�4�%�VJ�F��{���TO��.ȅ��J�NȎs�B
 M�g5��%�M_Y/�^�¹�e���3�xF����F�P� b��Z��+�q�r��=8��A�̙�;�y�>�����G_nm�,��j��t;��!����m^6N���*Ƈw;ո�����N�$�Ƣ�/몍N�������d�����.|d�X�B�����~Q�Xl=O�@��²a��Ȃ�9�(Y�G�E�j����oߙ�(ml���d����H���x�a�*r8��k��=�T��:���d�����`�W�\�e0;�ߘ�O����d�C=3�`g������{s�b�Y>�fW@aZ�]�^�Y/�^�¹�e���3S��T,c�z����Pq4^y@�c;҉��*��?$�B��u|����$�1X;��|B�'��|b�o�alֶ5mL^��a�@�nb:�N�NL�^	��a.�?�d���&��v�<��$�&�̞Y�&T�ͪ͌��LQ�qRN�-��º�Sr��nt��!�T�.��B�
/Sq�d��l����v�}�T�b����1��a"�!���ʵ�����dH�L�p��HM�ex�*aE�@[�_zβr�j5�{�0����%���p7���!���睋2'B�I��g?	��o�dEr�+��#ȕ�B N��r*�UӇ��ɋ� ��X�D
CvK}D�B��U������z*��['D�C�k�a�	�+4D@>�ܖ�4���D�gZ�w�q9+t�}t���3�l��d��JXl'�&�P�2�PUг�|<�D�$0����}�b�;�N�cP�`pJ����
@����=7�}|��	��a-6�Da�_.���%�줝v)��ɛ�?ө�Kf
�fWxxܤ�]
���b�v���V�i�;�H���o�4�= w
��ݔ��������@/��r �,fc�i���+J�2�f�;�>)�ӔuP��N�
�!���i��ċ�!-M�O��~��D�$0�y�R�QY`�CgD�|A�$����@/��r ��%�z�J��M:cD���Ȇb�L�($Z�u��΄x�g��	��S8�M�����vg����PTse��ͳ[�%�z�J��K�F�ش���R�t����ʵ������v�Z鎬�������(�����?�cc��L=X�� �-M�O��~�r�^�#v��.ȅ��J���B�:����}7�������\�2���.Z��'#P�j2E�?��˓#���l����d���=|%��v��3t���=�4�04�jfrw�&�z<a�4�ڈti@`:v�eQ۞h�G��#@�h�R*E���&�Ut�\�@�\����Ԍ��Ǐ�c���w�I�7z��,fqJ�jK�o[���[�2ٿ�VS`��@/��r ��%�z�J���,2�C�����d���Ą�Ĺ�,7�cL���	Ǹ�y85��n���d����P�ħN�g�c�`C��׍�߃��:����k������'#5��!�q�2��Kk:)���2�z�X
3kZ�T۳�͕���]�UQ��D�gZ�w�q9+t�}�xȀ��D׏�����Mp�-a�D͢q��`�L�5ߧE4��rw�&�z<a��N� ��靤�}O��ܐ�}�q���C�(�o�>�������7Ǧ���0+C��q��®��f�;�>)�L�N��Ѯy=k�Rm����s
!����p�>�q�M�4����3Urj��[R�03��ګ@�_kn��
���t׭Ҵ��=���D����\O]��S����7��@���kJU�4{��F	<���Hn
V~$
�8�O��Ίѥ֤�g�꿁��Ȝxڣ9�$���>��o���/i�D�]
���b��c���f�;�>)�ӔuP��Ni��ċ�!-M�O��~�Ѩ�f?�R�Ԍ��Ǐ�c���w�I�7['D�C�k�a�	�+4D@��"n�Κ�PޟT��&��,otFng��	T��Kf
�fKr���їu�ǏX����S)�3=7�}|��	m [}�؏[b%Ɨ����������O6��G�ez��2���թ�~X���@&�>�a���j_���N�K����3ύ\0K��̖���i��"u���Ȇb�L�($Z�u��΄x�g��	��S8�>���r8j�g����PTse��ͳ[�%�z�J���,2�C���l�yi��L.bC��k�]��^LP6݃۷��%�z�J���zt��[�6ZVE���Xu���#P�j2E�?��˓#���)��]ӈ�$I��}D�&�jW� ��z=���x(�i��/Rn����k���# m>���^!� wٻKm�Xn�
c����^eJ7�q���gҽd6�Kf
�f� *�P����j�1>�+�9-�i"'���Xw�j�7��#�@(14~�����-/J�����Ut�\�T۳�͕��)��]ӈ��s+N����Y�J������Q����ۉy�T�i��qolωP�HS|�4�04�jfJ�1����ݾ-/�uu��ڿ׏�����M��ܐ�}�6߳v�F���'��*��tw:g�V|�hi��p�7��Z鎬�����R�LM��ħƿ�9c�1��8�h�� ����f�#�eM�f<�,=K�F~�?|�[_c9��*��OT��]S��SO,F=d�g4"<·��3��J��@���,��t+����� ��P�!���2��O�O�d��,U��2�>D�c�lQw�v�����zL͊�q����N�:�Pn������Y�
�b9���:&�>��s����ӓ��^hq��:0k�y��HzL͊�q���@F�4��d��X���n���m!iI�"�,�>E��<��z��}�Q2�+�Y��c���9������5	��]�!��s[RTP��0c�,�[`������
L'���Xw�j�7����2�K<3�,P�zh�g��U-�e�TL���Y.��, #3������ls^3����� Oag�qod�֓��)b��X �<�3եt��'�=E1�r,��>T�ѐJj���Y�{'%sgeߪ�{ ^�x~�(vi�t�c,�q�T�\ ��9O���t�6�my$�N���Uە���׎o�|�ug�W���]�!��	Ǹ�y85���4
B<�%鯅�N�*�[Z�u�ZY�����Ayv߆��S&ϊu�z��[cƉ��#�Tۡ0�bm����e��3��v�/Q,��x��3����Hhqu!���5�Nn���4L"�#W��xW�Kg!�h�����7�$�G�j/����X�e��}c���G��m\Ӓ�qܛ�	����(:��=�M��0�d�Sd��_�a���n�|Wg�|bVzN7	+`�9
EMܓ���;�e >���l�n�Zl��Ͳ�8�3
�{�-�>��t��ԱͽP�nT��Э��y�L*���8�^�.eO��q��S��;�(e)��v��=����'�$��u,��y�"���Չ-d��r�b+��/6!��Ei�gz�����n�|W;"V7��evwJ���&�o�\,9o$aϛ`!�A���
+,I�2Sj�	�$ɜ�\�۟�-?�d���&����{ԕ�h7�{`��������* -��ed.:E������ƄH����[��2����s�Z΃xI��o�.�����U��)��d��y5\a�L�WStԪ���l���d��JXl'�&�P�2�PUг�|<q܃NQq�Je��v��$����Ze?&)�5#ғD+���4Y!�`�(i3!�`�(i3�����L�	�=����k�\Dc}՟2R��I���f(7���	�M|Y�N\��
�M�f��d,(!�`�(i3RN�]�5'���j���J�1��j��G��9B �b�ϧ��T�G��9B v�qi�S������|���k���Ô��xl}�<�9�t�Z��P���<�=z��jbkAޚN��^�ۍ�t���Q��S�����̲T��k��I�N��	T�i�Z�&�$I��h\���p>T!�`�(i3!�`�(i3nTxꅗ�~Fa�6"{�s��l���g�8> �T� 288��������k��&�Z�ӺVpaUv���Q�O='�)�����)��yG�%���!j��gÁ�r���Gg�o�Ɵ����J�F�c��4� wx�����nδ���5C!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3+Xz�4�焑�6G4��3> հ�`�H<�b��oW<���>��Z{��3�����Q�r�yK�9��7�_���.":�!�`�(i3!�`�(i3�`�>'r�:�;�ࢄH��L�}�?�}�r�2�"��Тϫ��8��/�	�d�H�K!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�����L�	u]�MP��br6��ۻ 288����Se�9'�ʺ&�Z�Ӻ�;�N�cP��8��	͂'�)�����?�}�r�2%���!j�Q.�U*Y�!�`�(i3!�`�(i3rz��G�x�����nδ���5CA
��z(����-@���m-NJ�*�#��d~�/�v�)�BҺ�)�|�$)#�o���!�`�(i3!�`�(i3!�`�(i3!�`�(i3�%_Z�ք{q��#�i+����Ó�d+st�I6�3> հ�`�H<�b�uu��N�B�>��Z{��A
��z(�k�dF�~"!�`�(i3!�`�(i3!�`�(i3!�`�(i3����k��J�Z���>H��L�}Q.�U*Y��"��Тϫ��8��/�R��\ !�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�����L�	�U��x]�i�A�Q�8�� 288����Z���u��&�Z�ӺA
��z(���I���'�)�����Q.�U*Y�!�`�(i3!�`�(i3!�`�(i3!�`�(i3rz��G�;����A=&�������!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3+Xz�4��W�i��8t�3> հ�`�H<�b���ˢYۋ!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�`�>'r�:�;�ࢄH��L�}���V�Ĩ"��Тϫ��8��/�I�$�jܲ!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�����L�	u]�MP��br6��ۻ 288���ɚ�ؘ�_�&�Z�Ӻk��=����8��	͂'�)��������V��%���!j��;t�b��!�`�(i3!�`�(i3rz��G�x�����nδ���5CA
��z(��������m-NJ�*�p�������v�)�BҺ�)�|�$��Y�c�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�%_Z�ք{q��#�i+����Ó�%���d��G�3> հ�`�H<�b��<��K��w�>��Z{��A
��z(�����VJ��!�`�(i3!�`�(i3!�`�(i3!�`�(i3����k��J�Z���>H��L�}�;t�b���"��Тϫ��8��/�kB��n&!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�����L�	�U��x]�i�A�Q�8�� 288����pq���:�&�Z�ӺA
��z(���qJ��
'�)�����;t�b��!�`�(i3!�`�(i3!�`�(i3!�`�(i3rz��G�;����A=&��B�Q�p׏�����M��ܐ�}����J���+)���܄���9<�f퀔������	-$ߔ���e�cN�\V����{�I�e5:�L��L�q���<�{�!���"�o��]gKl۞h�G��!�REK9�ӧK�or��	P�����9D�:��F�ā��O�q�V���p����z��-����C�;��GN�Y�,P�zh�g��U-�ea�}x2��VU�簦-�b�+�