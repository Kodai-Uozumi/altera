library verilog;
use verilog.vl_types.all;
entity \FILTER\ is
    port(
        \Y\             : out    vl_logic;
        \IN1\           : in     vl_logic
    );
end \FILTER\;
