library verilog;
use verilog.vl_types.all;
entity \TRIBUF\ is
    port(
        \Y\             : out    vl_logic;
        \IN1\           : in     vl_logic;
        \OE\            : in     vl_logic
    );
end \TRIBUF\;
